
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_unsigned.all;

entity top is 
end top;

architecture top of top is

---- Component declarations -----

component branch_unit
  port (
       A : in STD_LOGIC_VECTOR(127 downto 0);
       I16 : in STD_LOGIC_VECTOR(15 downto 0);
       PC : in STD_LOGIC_VECTOR(31 downto 0);
       T : in STD_LOGIC_VECTOR(127 downto 0);
       op_sel : in STD_LOGIC_VECTOR(2 downto 0);
       Result : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;
component byte_unit
  port (
       A : in STD_LOGIC_VECTOR(127 downto 0);
       B : in STD_LOGIC_VECTOR(127 downto 0);
       op_sel : in STD_LOGIC_VECTOR(1 downto 0);
       Result : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;
component even_pipe_reg
  port (
       Latency_d : in STD_LOGIC_VECTOR(2 downto 0);
       RegWr_d : in STD_LOGIC;
       RegdDst_d : in STD_LOGIC_VECTOR(6 downto 0);
       Result_d : in STD_LOGIC_VECTOR(127 downto 0);
       Unit_d : in STD_LOGIC_VECTOR(2 downto 0);
       clk : in STD_LOGIC;
       Latency_q : out STD_LOGIC_VECTOR(2 downto 0);
       RegWr_q : out STD_LOGIC;
       RegdDst_q : out STD_LOGIC_VECTOR(6 downto 0);
       Result_q : out STD_LOGIC_VECTOR(127 downto 0);
       Unit_q : out STD_LOGIC_VECTOR(2 downto 0)
  );
end component;
component forwarding_unit
  port (
       A_reg : in STD_LOGIC_VECTOR(127 downto 0);
       B_reg : in STD_LOGIC_VECTOR(127 downto 0);
       C_reg : in STD_LOGIC_VECTOR(127 downto 0);
       D_reg : in STD_LOGIC_VECTOR(127 downto 0);
       E_reg : in STD_LOGIC_VECTOR(127 downto 0);
       F_reg : in STD_LOGIC_VECTOR(127 downto 0);
       RA : in STD_LOGIC_VECTOR(6 downto 0);
       RB : in STD_LOGIC_VECTOR(6 downto 0);
       RC : in STD_LOGIC_VECTOR(6 downto 0);
       RD : in STD_LOGIC_VECTOR(6 downto 0);
       RE : in STD_LOGIC_VECTOR(6 downto 0);
       RF : in STD_LOGIC_VECTOR(6 downto 0);
       even1_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       even1_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       even1_RegWr : in STD_LOGIC;
       even1_Result : in STD_LOGIC_VECTOR(127 downto 0);
       even2_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       even2_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       even2_RegWr : in STD_LOGIC;
       even2_Result : in STD_LOGIC_VECTOR(127 downto 0);
       even3_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       even3_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       even3_RegWr : in STD_LOGIC;
       even3_Result : in STD_LOGIC_VECTOR(127 downto 0);
       even4_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       even4_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       even4_RegWr : in STD_LOGIC;
       even4_Result : in STD_LOGIC_VECTOR(127 downto 0);
       even5_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       even5_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       even5_RegWr : in STD_LOGIC;
       even5_Result : in STD_LOGIC_VECTOR(127 downto 0);
       even6_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       even6_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       even6_RegWr : in STD_LOGIC;
       even6_Result : in STD_LOGIC_VECTOR(127 downto 0);
       even7_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       even7_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       even7_RegWr : in STD_LOGIC;
       even7_Result : in STD_LOGIC_VECTOR(127 downto 0);
       odd1_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       odd1_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       odd1_RegWr : in STD_LOGIC;
       odd1_Result : in STD_LOGIC_VECTOR(127 downto 0);
       odd2_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       odd2_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       odd2_RegWr : in STD_LOGIC;
       odd2_Result : in STD_LOGIC_VECTOR(127 downto 0);
       odd3_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       odd3_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       odd3_RegWr : in STD_LOGIC;
       odd3_Result : in STD_LOGIC_VECTOR(127 downto 0);
       odd4_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       odd4_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       odd4_RegWr : in STD_LOGIC;
       odd4_Result : in STD_LOGIC_VECTOR(127 downto 0);
       odd5_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       odd5_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       odd5_RegWr : in STD_LOGIC;
       odd5_Result : in STD_LOGIC_VECTOR(127 downto 0);
       odd6_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       odd6_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       odd6_RegWr : in STD_LOGIC;
       odd6_Result : in STD_LOGIC_VECTOR(127 downto 0);
       odd7_Latency : in STD_LOGIC_VECTOR(2 downto 0);
       odd7_RegDst : in STD_LOGIC_VECTOR(6 downto 0);
       odd7_RegWr : in STD_LOGIC;
       odd7_Result : in STD_LOGIC_VECTOR(127 downto 0);
       A : out STD_LOGIC_VECTOR(127 downto 0);
       B : out STD_LOGIC_VECTOR(127 downto 0);
       C : out STD_LOGIC_VECTOR(127 downto 0);
       D : out STD_LOGIC_VECTOR(127 downto 0);
       E : out STD_LOGIC_VECTOR(127 downto 0);
       F : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;
component local_store_unit
  port (
       A : in STD_LOGIC_VECTOR(127 downto 0);
       B : in STD_LOGIC_VECTOR(127 downto 0);
       I10 : in STD_LOGIC_VECTOR(9 downto 0);
       I16 : in STD_LOGIC_VECTOR(15 downto 0);
       T : in STD_LOGIC_VECTOR(127 downto 0);
       clk : in STD_LOGIC;
       op_sel : in STD_LOGIC_VECTOR(2 downto 0);
       Result : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;
component odd_pipe_reg
  port (
       Branch_d : in STD_LOGIC;
       Latency_d : in STD_LOGIC_VECTOR(2 downto 0);
       RegWr_d : in STD_LOGIC;
       RegdDst_d : in STD_LOGIC_VECTOR(6 downto 0);
       Result_d : in STD_LOGIC_VECTOR(127 downto 0);
       Unit_d : in STD_LOGIC_VECTOR(2 downto 0);
       clk : in STD_LOGIC;
       Branch_q : out STD_LOGIC;
       Latency_q : out STD_LOGIC_VECTOR(2 downto 0);
       RegWr_q : out STD_LOGIC;
       RegdDst_q : out STD_LOGIC_VECTOR(6 downto 0);
       Result_q : out STD_LOGIC_VECTOR(127 downto 0);
       Unit_q : out STD_LOGIC_VECTOR(2 downto 0)
  );
end component;
component permute_unit
  port (
       A : in STD_LOGIC_VECTOR(127 downto 0);
       op_sel : in STD_LOGIC_VECTOR(1 downto 0);
       Result : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;
component register_file
  port (
       A_rd_addr : in STD_LOGIC_VECTOR(6 downto 0);
       A_wr_addr : in STD_LOGIC_VECTOR(6 downto 0);
       A_wr_data : in STD_LOGIC_VECTOR(127 downto 0);
       A_wr_en : in STD_LOGIC;
       B_rd_addr : in STD_LOGIC_VECTOR(6 downto 0);
       B_wr_addr : in STD_LOGIC_VECTOR(6 downto 0);
       B_wr_data : in STD_LOGIC_VECTOR(127 downto 0);
       B_wr_en : in STD_LOGIC;
       C_rd_addr : in STD_LOGIC_VECTOR(6 downto 0);
       D_rd_addr : in STD_LOGIC_VECTOR(6 downto 0);
       E_rd_addr : in STD_LOGIC_VECTOR(6 downto 0);
       F_rd_addr : in STD_LOGIC_VECTOR(6 downto 0);
       clk : in STD_LOGIC;
       A_rd_data : out STD_LOGIC_VECTOR(127 downto 0);
       B_rd_data : out STD_LOGIC_VECTOR(127 downto 0);
       C_rd_data : out STD_LOGIC_VECTOR(127 downto 0);
       D_rd_data : out STD_LOGIC_VECTOR(127 downto 0);
       E_rd_data : out STD_LOGIC_VECTOR(127 downto 0);
       F_rd_data : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;
component simple_fixed_unit1
  port (
       A : in STD_LOGIC_VECTOR(127 downto 0);
       B : in STD_LOGIC_VECTOR(127 downto 0);
       I10 : in STD_LOGIC_VECTOR(9 downto 0);
       I16 : in STD_LOGIC_VECTOR(15 downto 0);
       I18 : in STD_LOGIC_VECTOR(17 downto 0);
       op_sel : in STD_LOGIC_VECTOR(4 downto 0);
       Result : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;
component simple_fixed_unit2
  port (
       A : in STD_LOGIC_VECTOR(127 downto 0);
       B : in STD_LOGIC_VECTOR(127 downto 0);
       I7 : in STD_LOGIC_VECTOR(6 downto 0);
       op_sel : in STD_LOGIC_VECTOR(2 downto 0);
       Result : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;
component single_precision_unit
  port (
       A : in STD_LOGIC_VECTOR(127 downto 0);
       B : in STD_LOGIC_VECTOR(127 downto 0);
       C : in STD_LOGIC_VECTOR(127 downto 0);
       I10 : in STD_LOGIC_VECTOR(9 downto 0);
       I8 : in STD_LOGIC_VECTOR(7 downto 0);
       op_sel : in STD_LOGIC_VECTOR(3 downto 0);
       Result : out STD_LOGIC_VECTOR(127 downto 0)
  );
end component;

----     Constants     -----
constant DANGLING_INPUT_CONSTANT : STD_LOGIC := 'Z';

---- Signal declarations used on the diagram ----

signal A_wr_en : STD_LOGIC;
signal B_wr_en : STD_LOGIC;
signal NET1703 : STD_LOGIC;
signal NET1711 : STD_LOGIC;
signal NET600 : STD_LOGIC;
signal A_wr_addr : STD_LOGIC_VECTOR(6 downto 0);
signal A_wr_data : STD_LOGIC_VECTOR(127 downto 0);
signal BUS1695 : STD_LOGIC_VECTOR(6 downto 0);
signal BUS1719 : STD_LOGIC_VECTOR(2 downto 0);
signal BUS1766 : STD_LOGIC_VECTOR(6 downto 0);
signal BUS1770 : STD_LOGIC_VECTOR(6 downto 0);
signal BUS1774 : STD_LOGIC_VECTOR(6 downto 0);
signal BUS1778 : STD_LOGIC_VECTOR(6 downto 0);
signal BUS1782 : STD_LOGIC_VECTOR(6 downto 0);
signal BUS1786 : STD_LOGIC_VECTOR(7 downto 0);
signal BUS1961 : STD_LOGIC_VECTOR(2 downto 0);
signal BUS2032 : STD_LOGIC_VECTOR(7 downto 0);
signal BUS209 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS245 : STD_LOGIC_VECTOR(7 downto 0);
signal BUS297 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS328 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS331 : STD_LOGIC_VECTOR(9 downto 0);
signal BUS608 : STD_LOGIC_VECTOR(6 downto 0);
signal BUS616 : STD_LOGIC_VECTOR(1 downto 0);
signal BUS620 : STD_LOGIC_VECTOR(3 downto 0);
signal BUS624 : STD_LOGIC_VECTOR(2 downto 0);
signal BUS628 : STD_LOGIC_VECTOR(4 downto 0);
signal BUS632 : STD_LOGIC_VECTOR(15 downto 0);
signal BUS636 : STD_LOGIC_VECTOR(17 downto 0);
signal BUS640 : STD_LOGIC_VECTOR(6 downto 0);
signal BUS644 : STD_LOGIC_VECTOR(7 downto 0);
signal BUS648 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS670 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS678 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS686 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS694 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS709 : STD_LOGIC_VECTOR(2 downto 0);
signal BUS725 : STD_LOGIC_VECTOR(1 downto 0);
signal BUS733 : STD_LOGIC_VECTOR(2 downto 0);
signal BUS741 : STD_LOGIC_VECTOR(31 downto 0);
signal BUS751 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS758 : STD_LOGIC_VECTOR(2 downto 0);
signal BUS762 : STD_LOGIC_VECTOR(9 downto 0);
signal BUS772 : STD_LOGIC_VECTOR(15 downto 0);
signal BUS779 : STD_LOGIC_VECTOR(127 downto 0);
signal BUS789 : STD_LOGIC_VECTOR(127 downto 0);
signal B_wr_addr : STD_LOGIC_VECTOR(6 downto 0);
signal B_wr_data : STD_LOGIC_VECTOR(127 downto 0);

---- Declaration for Dangling input ----
signal Dangling_Input_Signal : STD_LOGIC;

---- Declarations for Dangling outputs ----
signal DANGLING_U33_Result_119 : STD_LOGIC;
signal DANGLING_U33_Result_118 : STD_LOGIC;
signal DANGLING_U33_Result_117 : STD_LOGIC;
signal DANGLING_U33_Result_116 : STD_LOGIC;
signal DANGLING_U33_Result_115 : STD_LOGIC;
signal DANGLING_U33_Result_114 : STD_LOGIC;
signal DANGLING_U33_Result_113 : STD_LOGIC;
signal DANGLING_U33_Result_112 : STD_LOGIC;
signal DANGLING_U33_Result_111 : STD_LOGIC;
signal DANGLING_U33_Result_110 : STD_LOGIC;
signal DANGLING_U33_Result_109 : STD_LOGIC;
signal DANGLING_U33_Result_108 : STD_LOGIC;
signal DANGLING_U33_Result_107 : STD_LOGIC;
signal DANGLING_U33_Result_106 : STD_LOGIC;
signal DANGLING_U33_Result_105 : STD_LOGIC;
signal DANGLING_U33_Result_104 : STD_LOGIC;
signal DANGLING_U33_Result_103 : STD_LOGIC;
signal DANGLING_U33_Result_102 : STD_LOGIC;
signal DANGLING_U33_Result_101 : STD_LOGIC;
signal DANGLING_U33_Result_100 : STD_LOGIC;
signal DANGLING_U33_Result_99 : STD_LOGIC;
signal DANGLING_U33_Result_98 : STD_LOGIC;
signal DANGLING_U33_Result_97 : STD_LOGIC;
signal DANGLING_U33_Result_96 : STD_LOGIC;
signal DANGLING_U33_Result_95 : STD_LOGIC;
signal DANGLING_U33_Result_94 : STD_LOGIC;
signal DANGLING_U33_Result_93 : STD_LOGIC;
signal DANGLING_U33_Result_92 : STD_LOGIC;
signal DANGLING_U33_Result_91 : STD_LOGIC;
signal DANGLING_U33_Result_90 : STD_LOGIC;
signal DANGLING_U33_Result_89 : STD_LOGIC;
signal DANGLING_U33_Result_88 : STD_LOGIC;
signal DANGLING_U33_Result_87 : STD_LOGIC;
signal DANGLING_U33_Result_86 : STD_LOGIC;
signal DANGLING_U33_Result_85 : STD_LOGIC;
signal DANGLING_U33_Result_84 : STD_LOGIC;
signal DANGLING_U33_Result_83 : STD_LOGIC;
signal DANGLING_U33_Result_82 : STD_LOGIC;
signal DANGLING_U33_Result_81 : STD_LOGIC;
signal DANGLING_U33_Result_80 : STD_LOGIC;
signal DANGLING_U33_Result_79 : STD_LOGIC;
signal DANGLING_U33_Result_78 : STD_LOGIC;
signal DANGLING_U33_Result_77 : STD_LOGIC;
signal DANGLING_U33_Result_76 : STD_LOGIC;
signal DANGLING_U33_Result_75 : STD_LOGIC;
signal DANGLING_U33_Result_74 : STD_LOGIC;
signal DANGLING_U33_Result_73 : STD_LOGIC;
signal DANGLING_U33_Result_72 : STD_LOGIC;
signal DANGLING_U33_Result_71 : STD_LOGIC;
signal DANGLING_U33_Result_70 : STD_LOGIC;
signal DANGLING_U33_Result_69 : STD_LOGIC;
signal DANGLING_U33_Result_68 : STD_LOGIC;
signal DANGLING_U33_Result_67 : STD_LOGIC;
signal DANGLING_U33_Result_66 : STD_LOGIC;
signal DANGLING_U33_Result_65 : STD_LOGIC;
signal DANGLING_U33_Result_64 : STD_LOGIC;
signal DANGLING_U33_Result_63 : STD_LOGIC;
signal DANGLING_U33_Result_62 : STD_LOGIC;
signal DANGLING_U33_Result_61 : STD_LOGIC;
signal DANGLING_U33_Result_60 : STD_LOGIC;
signal DANGLING_U33_Result_59 : STD_LOGIC;
signal DANGLING_U33_Result_58 : STD_LOGIC;
signal DANGLING_U33_Result_57 : STD_LOGIC;
signal DANGLING_U33_Result_56 : STD_LOGIC;
signal DANGLING_U33_Result_55 : STD_LOGIC;
signal DANGLING_U33_Result_54 : STD_LOGIC;
signal DANGLING_U33_Result_53 : STD_LOGIC;
signal DANGLING_U33_Result_52 : STD_LOGIC;
signal DANGLING_U33_Result_51 : STD_LOGIC;
signal DANGLING_U33_Result_50 : STD_LOGIC;
signal DANGLING_U33_Result_49 : STD_LOGIC;
signal DANGLING_U33_Result_48 : STD_LOGIC;
signal DANGLING_U33_Result_47 : STD_LOGIC;
signal DANGLING_U33_Result_46 : STD_LOGIC;
signal DANGLING_U33_Result_45 : STD_LOGIC;
signal DANGLING_U33_Result_44 : STD_LOGIC;
signal DANGLING_U33_Result_43 : STD_LOGIC;
signal DANGLING_U33_Result_42 : STD_LOGIC;
signal DANGLING_U33_Result_41 : STD_LOGIC;
signal DANGLING_U33_Result_40 : STD_LOGIC;
signal DANGLING_U33_Result_39 : STD_LOGIC;
signal DANGLING_U33_Result_38 : STD_LOGIC;
signal DANGLING_U33_Result_37 : STD_LOGIC;
signal DANGLING_U33_Result_36 : STD_LOGIC;
signal DANGLING_U33_Result_35 : STD_LOGIC;
signal DANGLING_U33_Result_34 : STD_LOGIC;
signal DANGLING_U33_Result_33 : STD_LOGIC;
signal DANGLING_U33_Result_32 : STD_LOGIC;
signal DANGLING_U33_Result_31 : STD_LOGIC;
signal DANGLING_U33_Result_30 : STD_LOGIC;
signal DANGLING_U33_Result_29 : STD_LOGIC;
signal DANGLING_U33_Result_28 : STD_LOGIC;
signal DANGLING_U33_Result_27 : STD_LOGIC;
signal DANGLING_U33_Result_26 : STD_LOGIC;
signal DANGLING_U33_Result_25 : STD_LOGIC;
signal DANGLING_U33_Result_24 : STD_LOGIC;
signal DANGLING_U33_Result_23 : STD_LOGIC;
signal DANGLING_U33_Result_22 : STD_LOGIC;
signal DANGLING_U33_Result_21 : STD_LOGIC;
signal DANGLING_U33_Result_20 : STD_LOGIC;
signal DANGLING_U33_Result_19 : STD_LOGIC;
signal DANGLING_U33_Result_18 : STD_LOGIC;
signal DANGLING_U33_Result_17 : STD_LOGIC;
signal DANGLING_U33_Result_16 : STD_LOGIC;
signal DANGLING_U33_Result_15 : STD_LOGIC;
signal DANGLING_U33_Result_14 : STD_LOGIC;
signal DANGLING_U33_Result_13 : STD_LOGIC;
signal DANGLING_U33_Result_12 : STD_LOGIC;
signal DANGLING_U33_Result_11 : STD_LOGIC;
signal DANGLING_U33_Result_10 : STD_LOGIC;
signal DANGLING_U33_Result_9 : STD_LOGIC;
signal DANGLING_U33_Result_8 : STD_LOGIC;
signal DANGLING_U33_Result_7 : STD_LOGIC;
signal DANGLING_U33_Result_6 : STD_LOGIC;
signal DANGLING_U33_Result_5 : STD_LOGIC;
signal DANGLING_U33_Result_4 : STD_LOGIC;
signal DANGLING_U33_Result_3 : STD_LOGIC;
signal DANGLING_U33_Result_2 : STD_LOGIC;
signal DANGLING_U33_Result_1 : STD_LOGIC;
signal DANGLING_U33_Result_0 : STD_LOGIC;
signal DANGLING_U34_Result_119 : STD_LOGIC;
signal DANGLING_U34_Result_118 : STD_LOGIC;
signal DANGLING_U34_Result_117 : STD_LOGIC;
signal DANGLING_U34_Result_116 : STD_LOGIC;
signal DANGLING_U34_Result_115 : STD_LOGIC;
signal DANGLING_U34_Result_114 : STD_LOGIC;
signal DANGLING_U34_Result_113 : STD_LOGIC;
signal DANGLING_U34_Result_112 : STD_LOGIC;
signal DANGLING_U34_Result_111 : STD_LOGIC;
signal DANGLING_U34_Result_110 : STD_LOGIC;
signal DANGLING_U34_Result_109 : STD_LOGIC;
signal DANGLING_U34_Result_108 : STD_LOGIC;
signal DANGLING_U34_Result_107 : STD_LOGIC;
signal DANGLING_U34_Result_106 : STD_LOGIC;
signal DANGLING_U34_Result_105 : STD_LOGIC;
signal DANGLING_U34_Result_104 : STD_LOGIC;
signal DANGLING_U34_Result_103 : STD_LOGIC;
signal DANGLING_U34_Result_102 : STD_LOGIC;
signal DANGLING_U34_Result_101 : STD_LOGIC;
signal DANGLING_U34_Result_100 : STD_LOGIC;
signal DANGLING_U34_Result_99 : STD_LOGIC;
signal DANGLING_U34_Result_98 : STD_LOGIC;
signal DANGLING_U34_Result_97 : STD_LOGIC;
signal DANGLING_U34_Result_96 : STD_LOGIC;
signal DANGLING_U34_Result_95 : STD_LOGIC;
signal DANGLING_U34_Result_94 : STD_LOGIC;
signal DANGLING_U34_Result_93 : STD_LOGIC;
signal DANGLING_U34_Result_92 : STD_LOGIC;
signal DANGLING_U34_Result_91 : STD_LOGIC;
signal DANGLING_U34_Result_90 : STD_LOGIC;
signal DANGLING_U34_Result_89 : STD_LOGIC;
signal DANGLING_U34_Result_88 : STD_LOGIC;
signal DANGLING_U34_Result_87 : STD_LOGIC;
signal DANGLING_U34_Result_86 : STD_LOGIC;
signal DANGLING_U34_Result_85 : STD_LOGIC;
signal DANGLING_U34_Result_84 : STD_LOGIC;
signal DANGLING_U34_Result_83 : STD_LOGIC;
signal DANGLING_U34_Result_82 : STD_LOGIC;
signal DANGLING_U34_Result_81 : STD_LOGIC;
signal DANGLING_U34_Result_80 : STD_LOGIC;
signal DANGLING_U34_Result_79 : STD_LOGIC;
signal DANGLING_U34_Result_78 : STD_LOGIC;
signal DANGLING_U34_Result_77 : STD_LOGIC;
signal DANGLING_U34_Result_76 : STD_LOGIC;
signal DANGLING_U34_Result_75 : STD_LOGIC;
signal DANGLING_U34_Result_74 : STD_LOGIC;
signal DANGLING_U34_Result_73 : STD_LOGIC;
signal DANGLING_U34_Result_72 : STD_LOGIC;
signal DANGLING_U34_Result_71 : STD_LOGIC;
signal DANGLING_U34_Result_70 : STD_LOGIC;
signal DANGLING_U34_Result_69 : STD_LOGIC;
signal DANGLING_U34_Result_68 : STD_LOGIC;
signal DANGLING_U34_Result_67 : STD_LOGIC;
signal DANGLING_U34_Result_66 : STD_LOGIC;
signal DANGLING_U34_Result_65 : STD_LOGIC;
signal DANGLING_U34_Result_64 : STD_LOGIC;
signal DANGLING_U34_Result_63 : STD_LOGIC;
signal DANGLING_U34_Result_62 : STD_LOGIC;
signal DANGLING_U34_Result_61 : STD_LOGIC;
signal DANGLING_U34_Result_60 : STD_LOGIC;
signal DANGLING_U34_Result_59 : STD_LOGIC;
signal DANGLING_U34_Result_58 : STD_LOGIC;
signal DANGLING_U34_Result_57 : STD_LOGIC;
signal DANGLING_U34_Result_56 : STD_LOGIC;
signal DANGLING_U34_Result_55 : STD_LOGIC;
signal DANGLING_U34_Result_54 : STD_LOGIC;
signal DANGLING_U34_Result_53 : STD_LOGIC;
signal DANGLING_U34_Result_52 : STD_LOGIC;
signal DANGLING_U34_Result_51 : STD_LOGIC;
signal DANGLING_U34_Result_50 : STD_LOGIC;
signal DANGLING_U34_Result_49 : STD_LOGIC;
signal DANGLING_U34_Result_48 : STD_LOGIC;
signal DANGLING_U34_Result_47 : STD_LOGIC;
signal DANGLING_U34_Result_46 : STD_LOGIC;
signal DANGLING_U34_Result_45 : STD_LOGIC;
signal DANGLING_U34_Result_44 : STD_LOGIC;
signal DANGLING_U34_Result_43 : STD_LOGIC;
signal DANGLING_U34_Result_42 : STD_LOGIC;
signal DANGLING_U34_Result_41 : STD_LOGIC;
signal DANGLING_U34_Result_40 : STD_LOGIC;
signal DANGLING_U34_Result_39 : STD_LOGIC;
signal DANGLING_U34_Result_38 : STD_LOGIC;
signal DANGLING_U34_Result_37 : STD_LOGIC;
signal DANGLING_U34_Result_36 : STD_LOGIC;
signal DANGLING_U34_Result_35 : STD_LOGIC;
signal DANGLING_U34_Result_34 : STD_LOGIC;
signal DANGLING_U34_Result_33 : STD_LOGIC;
signal DANGLING_U34_Result_32 : STD_LOGIC;
signal DANGLING_U34_Result_31 : STD_LOGIC;
signal DANGLING_U34_Result_30 : STD_LOGIC;
signal DANGLING_U34_Result_29 : STD_LOGIC;
signal DANGLING_U34_Result_28 : STD_LOGIC;
signal DANGLING_U34_Result_27 : STD_LOGIC;
signal DANGLING_U34_Result_26 : STD_LOGIC;
signal DANGLING_U34_Result_25 : STD_LOGIC;
signal DANGLING_U34_Result_24 : STD_LOGIC;
signal DANGLING_U34_Result_23 : STD_LOGIC;
signal DANGLING_U34_Result_22 : STD_LOGIC;
signal DANGLING_U34_Result_21 : STD_LOGIC;
signal DANGLING_U34_Result_20 : STD_LOGIC;
signal DANGLING_U34_Result_19 : STD_LOGIC;
signal DANGLING_U34_Result_18 : STD_LOGIC;
signal DANGLING_U34_Result_17 : STD_LOGIC;
signal DANGLING_U34_Result_16 : STD_LOGIC;
signal DANGLING_U34_Result_15 : STD_LOGIC;
signal DANGLING_U34_Result_14 : STD_LOGIC;
signal DANGLING_U34_Result_13 : STD_LOGIC;
signal DANGLING_U34_Result_12 : STD_LOGIC;
signal DANGLING_U34_Result_11 : STD_LOGIC;
signal DANGLING_U34_Result_10 : STD_LOGIC;
signal DANGLING_U34_Result_9 : STD_LOGIC;
signal DANGLING_U34_Result_8 : STD_LOGIC;
signal DANGLING_U34_Result_7 : STD_LOGIC;
signal DANGLING_U34_Result_6 : STD_LOGIC;
signal DANGLING_U34_Result_5 : STD_LOGIC;
signal DANGLING_U34_Result_4 : STD_LOGIC;
signal DANGLING_U34_Result_3 : STD_LOGIC;
signal DANGLING_U34_Result_2 : STD_LOGIC;
signal DANGLING_U34_Result_1 : STD_LOGIC;
signal DANGLING_U34_Result_0 : STD_LOGIC;
signal DANGLING_U35_Result_119 : STD_LOGIC;
signal DANGLING_U35_Result_118 : STD_LOGIC;
signal DANGLING_U35_Result_117 : STD_LOGIC;
signal DANGLING_U35_Result_116 : STD_LOGIC;
signal DANGLING_U35_Result_115 : STD_LOGIC;
signal DANGLING_U35_Result_114 : STD_LOGIC;
signal DANGLING_U35_Result_113 : STD_LOGIC;
signal DANGLING_U35_Result_112 : STD_LOGIC;
signal DANGLING_U35_Result_111 : STD_LOGIC;
signal DANGLING_U35_Result_110 : STD_LOGIC;
signal DANGLING_U35_Result_109 : STD_LOGIC;
signal DANGLING_U35_Result_108 : STD_LOGIC;
signal DANGLING_U35_Result_107 : STD_LOGIC;
signal DANGLING_U35_Result_106 : STD_LOGIC;
signal DANGLING_U35_Result_105 : STD_LOGIC;
signal DANGLING_U35_Result_104 : STD_LOGIC;
signal DANGLING_U35_Result_103 : STD_LOGIC;
signal DANGLING_U35_Result_102 : STD_LOGIC;
signal DANGLING_U35_Result_101 : STD_LOGIC;
signal DANGLING_U35_Result_100 : STD_LOGIC;
signal DANGLING_U35_Result_99 : STD_LOGIC;
signal DANGLING_U35_Result_98 : STD_LOGIC;
signal DANGLING_U35_Result_97 : STD_LOGIC;
signal DANGLING_U35_Result_96 : STD_LOGIC;
signal DANGLING_U35_Result_95 : STD_LOGIC;
signal DANGLING_U35_Result_94 : STD_LOGIC;
signal DANGLING_U35_Result_93 : STD_LOGIC;
signal DANGLING_U35_Result_92 : STD_LOGIC;
signal DANGLING_U35_Result_91 : STD_LOGIC;
signal DANGLING_U35_Result_90 : STD_LOGIC;
signal DANGLING_U35_Result_89 : STD_LOGIC;
signal DANGLING_U35_Result_88 : STD_LOGIC;
signal DANGLING_U35_Result_87 : STD_LOGIC;
signal DANGLING_U35_Result_86 : STD_LOGIC;
signal DANGLING_U35_Result_85 : STD_LOGIC;
signal DANGLING_U35_Result_84 : STD_LOGIC;
signal DANGLING_U35_Result_83 : STD_LOGIC;
signal DANGLING_U35_Result_82 : STD_LOGIC;
signal DANGLING_U35_Result_81 : STD_LOGIC;
signal DANGLING_U35_Result_80 : STD_LOGIC;
signal DANGLING_U35_Result_79 : STD_LOGIC;
signal DANGLING_U35_Result_78 : STD_LOGIC;
signal DANGLING_U35_Result_77 : STD_LOGIC;
signal DANGLING_U35_Result_76 : STD_LOGIC;
signal DANGLING_U35_Result_75 : STD_LOGIC;
signal DANGLING_U35_Result_74 : STD_LOGIC;
signal DANGLING_U35_Result_73 : STD_LOGIC;
signal DANGLING_U35_Result_72 : STD_LOGIC;
signal DANGLING_U35_Result_71 : STD_LOGIC;
signal DANGLING_U35_Result_70 : STD_LOGIC;
signal DANGLING_U35_Result_69 : STD_LOGIC;
signal DANGLING_U35_Result_68 : STD_LOGIC;
signal DANGLING_U35_Result_67 : STD_LOGIC;
signal DANGLING_U35_Result_66 : STD_LOGIC;
signal DANGLING_U35_Result_65 : STD_LOGIC;
signal DANGLING_U35_Result_64 : STD_LOGIC;
signal DANGLING_U35_Result_63 : STD_LOGIC;
signal DANGLING_U35_Result_62 : STD_LOGIC;
signal DANGLING_U35_Result_61 : STD_LOGIC;
signal DANGLING_U35_Result_60 : STD_LOGIC;
signal DANGLING_U35_Result_59 : STD_LOGIC;
signal DANGLING_U35_Result_58 : STD_LOGIC;
signal DANGLING_U35_Result_57 : STD_LOGIC;
signal DANGLING_U35_Result_56 : STD_LOGIC;
signal DANGLING_U35_Result_55 : STD_LOGIC;
signal DANGLING_U35_Result_54 : STD_LOGIC;
signal DANGLING_U35_Result_53 : STD_LOGIC;
signal DANGLING_U35_Result_52 : STD_LOGIC;
signal DANGLING_U35_Result_51 : STD_LOGIC;
signal DANGLING_U35_Result_50 : STD_LOGIC;
signal DANGLING_U35_Result_49 : STD_LOGIC;
signal DANGLING_U35_Result_48 : STD_LOGIC;
signal DANGLING_U35_Result_47 : STD_LOGIC;
signal DANGLING_U35_Result_46 : STD_LOGIC;
signal DANGLING_U35_Result_45 : STD_LOGIC;
signal DANGLING_U35_Result_44 : STD_LOGIC;
signal DANGLING_U35_Result_43 : STD_LOGIC;
signal DANGLING_U35_Result_42 : STD_LOGIC;
signal DANGLING_U35_Result_41 : STD_LOGIC;
signal DANGLING_U35_Result_40 : STD_LOGIC;
signal DANGLING_U35_Result_39 : STD_LOGIC;
signal DANGLING_U35_Result_38 : STD_LOGIC;
signal DANGLING_U35_Result_37 : STD_LOGIC;
signal DANGLING_U35_Result_36 : STD_LOGIC;
signal DANGLING_U35_Result_35 : STD_LOGIC;
signal DANGLING_U35_Result_34 : STD_LOGIC;
signal DANGLING_U35_Result_33 : STD_LOGIC;
signal DANGLING_U35_Result_32 : STD_LOGIC;
signal DANGLING_U35_Result_31 : STD_LOGIC;
signal DANGLING_U35_Result_30 : STD_LOGIC;
signal DANGLING_U35_Result_29 : STD_LOGIC;
signal DANGLING_U35_Result_28 : STD_LOGIC;
signal DANGLING_U35_Result_27 : STD_LOGIC;
signal DANGLING_U35_Result_26 : STD_LOGIC;
signal DANGLING_U35_Result_25 : STD_LOGIC;
signal DANGLING_U35_Result_24 : STD_LOGIC;
signal DANGLING_U35_Result_23 : STD_LOGIC;
signal DANGLING_U35_Result_22 : STD_LOGIC;
signal DANGLING_U35_Result_21 : STD_LOGIC;
signal DANGLING_U35_Result_20 : STD_LOGIC;
signal DANGLING_U35_Result_19 : STD_LOGIC;
signal DANGLING_U35_Result_18 : STD_LOGIC;
signal DANGLING_U35_Result_17 : STD_LOGIC;
signal DANGLING_U35_Result_16 : STD_LOGIC;
signal DANGLING_U35_Result_15 : STD_LOGIC;
signal DANGLING_U35_Result_14 : STD_LOGIC;
signal DANGLING_U35_Result_13 : STD_LOGIC;
signal DANGLING_U35_Result_12 : STD_LOGIC;
signal DANGLING_U35_Result_11 : STD_LOGIC;
signal DANGLING_U35_Result_10 : STD_LOGIC;
signal DANGLING_U35_Result_9 : STD_LOGIC;
signal DANGLING_U35_Result_8 : STD_LOGIC;
signal DANGLING_U35_Result_7 : STD_LOGIC;
signal DANGLING_U35_Result_6 : STD_LOGIC;
signal DANGLING_U35_Result_5 : STD_LOGIC;
signal DANGLING_U35_Result_4 : STD_LOGIC;
signal DANGLING_U35_Result_3 : STD_LOGIC;
signal DANGLING_U35_Result_2 : STD_LOGIC;
signal DANGLING_U35_Result_1 : STD_LOGIC;
signal DANGLING_U35_Result_0 : STD_LOGIC;

begin

----  Component instantiations  ----

U33 : simple_fixed_unit1
  port map(
       A => BUS328,
       B => BUS297,
       I10 => BUS331,
       I16 => BUS632,
       I18 => BUS636,
       Result(0) => DANGLING_U33_Result_0,
       Result(1) => DANGLING_U33_Result_1,
       Result(2) => DANGLING_U33_Result_2,
       Result(3) => DANGLING_U33_Result_3,
       Result(4) => DANGLING_U33_Result_4,
       Result(5) => DANGLING_U33_Result_5,
       Result(6) => DANGLING_U33_Result_6,
       Result(7) => DANGLING_U33_Result_7,
       Result(8) => DANGLING_U33_Result_8,
       Result(9) => DANGLING_U33_Result_9,
       Result(10) => DANGLING_U33_Result_10,
       Result(11) => DANGLING_U33_Result_11,
       Result(12) => DANGLING_U33_Result_12,
       Result(13) => DANGLING_U33_Result_13,
       Result(14) => DANGLING_U33_Result_14,
       Result(15) => DANGLING_U33_Result_15,
       Result(16) => DANGLING_U33_Result_16,
       Result(17) => DANGLING_U33_Result_17,
       Result(18) => DANGLING_U33_Result_18,
       Result(19) => DANGLING_U33_Result_19,
       Result(20) => DANGLING_U33_Result_20,
       Result(21) => DANGLING_U33_Result_21,
       Result(22) => DANGLING_U33_Result_22,
       Result(23) => DANGLING_U33_Result_23,
       Result(24) => DANGLING_U33_Result_24,
       Result(25) => DANGLING_U33_Result_25,
       Result(26) => DANGLING_U33_Result_26,
       Result(27) => DANGLING_U33_Result_27,
       Result(28) => DANGLING_U33_Result_28,
       Result(29) => DANGLING_U33_Result_29,
       Result(30) => DANGLING_U33_Result_30,
       Result(31) => DANGLING_U33_Result_31,
       Result(32) => DANGLING_U33_Result_32,
       Result(33) => DANGLING_U33_Result_33,
       Result(34) => DANGLING_U33_Result_34,
       Result(35) => DANGLING_U33_Result_35,
       Result(36) => DANGLING_U33_Result_36,
       Result(37) => DANGLING_U33_Result_37,
       Result(38) => DANGLING_U33_Result_38,
       Result(39) => DANGLING_U33_Result_39,
       Result(40) => DANGLING_U33_Result_40,
       Result(41) => DANGLING_U33_Result_41,
       Result(42) => DANGLING_U33_Result_42,
       Result(43) => DANGLING_U33_Result_43,
       Result(44) => DANGLING_U33_Result_44,
       Result(45) => DANGLING_U33_Result_45,
       Result(46) => DANGLING_U33_Result_46,
       Result(47) => DANGLING_U33_Result_47,
       Result(48) => DANGLING_U33_Result_48,
       Result(49) => DANGLING_U33_Result_49,
       Result(50) => DANGLING_U33_Result_50,
       Result(51) => DANGLING_U33_Result_51,
       Result(52) => DANGLING_U33_Result_52,
       Result(53) => DANGLING_U33_Result_53,
       Result(54) => DANGLING_U33_Result_54,
       Result(55) => DANGLING_U33_Result_55,
       Result(56) => DANGLING_U33_Result_56,
       Result(57) => DANGLING_U33_Result_57,
       Result(58) => DANGLING_U33_Result_58,
       Result(59) => DANGLING_U33_Result_59,
       Result(60) => DANGLING_U33_Result_60,
       Result(61) => DANGLING_U33_Result_61,
       Result(62) => DANGLING_U33_Result_62,
       Result(63) => DANGLING_U33_Result_63,
       Result(64) => DANGLING_U33_Result_64,
       Result(65) => DANGLING_U33_Result_65,
       Result(66) => DANGLING_U33_Result_66,
       Result(67) => DANGLING_U33_Result_67,
       Result(68) => DANGLING_U33_Result_68,
       Result(69) => DANGLING_U33_Result_69,
       Result(70) => DANGLING_U33_Result_70,
       Result(71) => DANGLING_U33_Result_71,
       Result(72) => DANGLING_U33_Result_72,
       Result(73) => DANGLING_U33_Result_73,
       Result(74) => DANGLING_U33_Result_74,
       Result(75) => DANGLING_U33_Result_75,
       Result(76) => DANGLING_U33_Result_76,
       Result(77) => DANGLING_U33_Result_77,
       Result(78) => DANGLING_U33_Result_78,
       Result(79) => DANGLING_U33_Result_79,
       Result(80) => DANGLING_U33_Result_80,
       Result(81) => DANGLING_U33_Result_81,
       Result(82) => DANGLING_U33_Result_82,
       Result(83) => DANGLING_U33_Result_83,
       Result(84) => DANGLING_U33_Result_84,
       Result(85) => DANGLING_U33_Result_85,
       Result(86) => DANGLING_U33_Result_86,
       Result(87) => DANGLING_U33_Result_87,
       Result(88) => DANGLING_U33_Result_88,
       Result(89) => DANGLING_U33_Result_89,
       Result(90) => DANGLING_U33_Result_90,
       Result(91) => DANGLING_U33_Result_91,
       Result(92) => DANGLING_U33_Result_92,
       Result(93) => DANGLING_U33_Result_93,
       Result(94) => DANGLING_U33_Result_94,
       Result(95) => DANGLING_U33_Result_95,
       Result(96) => DANGLING_U33_Result_96,
       Result(97) => DANGLING_U33_Result_97,
       Result(98) => DANGLING_U33_Result_98,
       Result(99) => DANGLING_U33_Result_99,
       Result(100) => DANGLING_U33_Result_100,
       Result(101) => DANGLING_U33_Result_101,
       Result(102) => DANGLING_U33_Result_102,
       Result(103) => DANGLING_U33_Result_103,
       Result(104) => DANGLING_U33_Result_104,
       Result(105) => DANGLING_U33_Result_105,
       Result(106) => DANGLING_U33_Result_106,
       Result(107) => DANGLING_U33_Result_107,
       Result(108) => DANGLING_U33_Result_108,
       Result(109) => DANGLING_U33_Result_109,
       Result(110) => DANGLING_U33_Result_110,
       Result(111) => DANGLING_U33_Result_111,
       Result(112) => DANGLING_U33_Result_112,
       Result(113) => DANGLING_U33_Result_113,
       Result(114) => DANGLING_U33_Result_114,
       Result(115) => DANGLING_U33_Result_115,
       Result(116) => DANGLING_U33_Result_116,
       Result(117) => DANGLING_U33_Result_117,
       Result(118) => DANGLING_U33_Result_118,
       Result(119) => DANGLING_U33_Result_119,
       Result(120) => BUS2032(0),
       Result(121) => BUS2032(1),
       Result(122) => BUS2032(2),
       Result(123) => BUS2032(3),
       Result(124) => BUS2032(4),
       Result(125) => BUS2032(5),
       Result(126) => BUS2032(6),
       Result(127) => BUS2032(7),
       op_sel => BUS628
  );

U34 : simple_fixed_unit2
  port map(
       A => BUS328,
       B => BUS297,
       I7 => BUS640,
       Result(0) => DANGLING_U34_Result_0,
       Result(1) => DANGLING_U34_Result_1,
       Result(2) => DANGLING_U34_Result_2,
       Result(3) => DANGLING_U34_Result_3,
       Result(4) => DANGLING_U34_Result_4,
       Result(5) => DANGLING_U34_Result_5,
       Result(6) => DANGLING_U34_Result_6,
       Result(7) => DANGLING_U34_Result_7,
       Result(8) => DANGLING_U34_Result_8,
       Result(9) => DANGLING_U34_Result_9,
       Result(10) => DANGLING_U34_Result_10,
       Result(11) => DANGLING_U34_Result_11,
       Result(12) => DANGLING_U34_Result_12,
       Result(13) => DANGLING_U34_Result_13,
       Result(14) => DANGLING_U34_Result_14,
       Result(15) => DANGLING_U34_Result_15,
       Result(16) => DANGLING_U34_Result_16,
       Result(17) => DANGLING_U34_Result_17,
       Result(18) => DANGLING_U34_Result_18,
       Result(19) => DANGLING_U34_Result_19,
       Result(20) => DANGLING_U34_Result_20,
       Result(21) => DANGLING_U34_Result_21,
       Result(22) => DANGLING_U34_Result_22,
       Result(23) => DANGLING_U34_Result_23,
       Result(24) => DANGLING_U34_Result_24,
       Result(25) => DANGLING_U34_Result_25,
       Result(26) => DANGLING_U34_Result_26,
       Result(27) => DANGLING_U34_Result_27,
       Result(28) => DANGLING_U34_Result_28,
       Result(29) => DANGLING_U34_Result_29,
       Result(30) => DANGLING_U34_Result_30,
       Result(31) => DANGLING_U34_Result_31,
       Result(32) => DANGLING_U34_Result_32,
       Result(33) => DANGLING_U34_Result_33,
       Result(34) => DANGLING_U34_Result_34,
       Result(35) => DANGLING_U34_Result_35,
       Result(36) => DANGLING_U34_Result_36,
       Result(37) => DANGLING_U34_Result_37,
       Result(38) => DANGLING_U34_Result_38,
       Result(39) => DANGLING_U34_Result_39,
       Result(40) => DANGLING_U34_Result_40,
       Result(41) => DANGLING_U34_Result_41,
       Result(42) => DANGLING_U34_Result_42,
       Result(43) => DANGLING_U34_Result_43,
       Result(44) => DANGLING_U34_Result_44,
       Result(45) => DANGLING_U34_Result_45,
       Result(46) => DANGLING_U34_Result_46,
       Result(47) => DANGLING_U34_Result_47,
       Result(48) => DANGLING_U34_Result_48,
       Result(49) => DANGLING_U34_Result_49,
       Result(50) => DANGLING_U34_Result_50,
       Result(51) => DANGLING_U34_Result_51,
       Result(52) => DANGLING_U34_Result_52,
       Result(53) => DANGLING_U34_Result_53,
       Result(54) => DANGLING_U34_Result_54,
       Result(55) => DANGLING_U34_Result_55,
       Result(56) => DANGLING_U34_Result_56,
       Result(57) => DANGLING_U34_Result_57,
       Result(58) => DANGLING_U34_Result_58,
       Result(59) => DANGLING_U34_Result_59,
       Result(60) => DANGLING_U34_Result_60,
       Result(61) => DANGLING_U34_Result_61,
       Result(62) => DANGLING_U34_Result_62,
       Result(63) => DANGLING_U34_Result_63,
       Result(64) => DANGLING_U34_Result_64,
       Result(65) => DANGLING_U34_Result_65,
       Result(66) => DANGLING_U34_Result_66,
       Result(67) => DANGLING_U34_Result_67,
       Result(68) => DANGLING_U34_Result_68,
       Result(69) => DANGLING_U34_Result_69,
       Result(70) => DANGLING_U34_Result_70,
       Result(71) => DANGLING_U34_Result_71,
       Result(72) => DANGLING_U34_Result_72,
       Result(73) => DANGLING_U34_Result_73,
       Result(74) => DANGLING_U34_Result_74,
       Result(75) => DANGLING_U34_Result_75,
       Result(76) => DANGLING_U34_Result_76,
       Result(77) => DANGLING_U34_Result_77,
       Result(78) => DANGLING_U34_Result_78,
       Result(79) => DANGLING_U34_Result_79,
       Result(80) => DANGLING_U34_Result_80,
       Result(81) => DANGLING_U34_Result_81,
       Result(82) => DANGLING_U34_Result_82,
       Result(83) => DANGLING_U34_Result_83,
       Result(84) => DANGLING_U34_Result_84,
       Result(85) => DANGLING_U34_Result_85,
       Result(86) => DANGLING_U34_Result_86,
       Result(87) => DANGLING_U34_Result_87,
       Result(88) => DANGLING_U34_Result_88,
       Result(89) => DANGLING_U34_Result_89,
       Result(90) => DANGLING_U34_Result_90,
       Result(91) => DANGLING_U34_Result_91,
       Result(92) => DANGLING_U34_Result_92,
       Result(93) => DANGLING_U34_Result_93,
       Result(94) => DANGLING_U34_Result_94,
       Result(95) => DANGLING_U34_Result_95,
       Result(96) => DANGLING_U34_Result_96,
       Result(97) => DANGLING_U34_Result_97,
       Result(98) => DANGLING_U34_Result_98,
       Result(99) => DANGLING_U34_Result_99,
       Result(100) => DANGLING_U34_Result_100,
       Result(101) => DANGLING_U34_Result_101,
       Result(102) => DANGLING_U34_Result_102,
       Result(103) => DANGLING_U34_Result_103,
       Result(104) => DANGLING_U34_Result_104,
       Result(105) => DANGLING_U34_Result_105,
       Result(106) => DANGLING_U34_Result_106,
       Result(107) => DANGLING_U34_Result_107,
       Result(108) => DANGLING_U34_Result_108,
       Result(109) => DANGLING_U34_Result_109,
       Result(110) => DANGLING_U34_Result_110,
       Result(111) => DANGLING_U34_Result_111,
       Result(112) => DANGLING_U34_Result_112,
       Result(113) => DANGLING_U34_Result_113,
       Result(114) => DANGLING_U34_Result_114,
       Result(115) => DANGLING_U34_Result_115,
       Result(116) => DANGLING_U34_Result_116,
       Result(117) => DANGLING_U34_Result_117,
       Result(118) => DANGLING_U34_Result_118,
       Result(119) => DANGLING_U34_Result_119,
       Result(120) => BUS2032(0),
       Result(121) => BUS2032(1),
       Result(122) => BUS2032(2),
       Result(123) => BUS2032(3),
       Result(124) => BUS2032(4),
       Result(125) => BUS2032(5),
       Result(126) => BUS2032(6),
       Result(127) => BUS2032(7),
       op_sel => BUS624
  );

U35 : single_precision_unit
  port map(
       A => BUS328,
       B => BUS297,
       C => BUS648,
       I10 => BUS331,
       I8 => BUS644,
       Result(0) => DANGLING_U35_Result_0,
       Result(1) => DANGLING_U35_Result_1,
       Result(2) => DANGLING_U35_Result_2,
       Result(3) => DANGLING_U35_Result_3,
       Result(4) => DANGLING_U35_Result_4,
       Result(5) => DANGLING_U35_Result_5,
       Result(6) => DANGLING_U35_Result_6,
       Result(7) => DANGLING_U35_Result_7,
       Result(8) => DANGLING_U35_Result_8,
       Result(9) => DANGLING_U35_Result_9,
       Result(10) => DANGLING_U35_Result_10,
       Result(11) => DANGLING_U35_Result_11,
       Result(12) => DANGLING_U35_Result_12,
       Result(13) => DANGLING_U35_Result_13,
       Result(14) => DANGLING_U35_Result_14,
       Result(15) => DANGLING_U35_Result_15,
       Result(16) => DANGLING_U35_Result_16,
       Result(17) => DANGLING_U35_Result_17,
       Result(18) => DANGLING_U35_Result_18,
       Result(19) => DANGLING_U35_Result_19,
       Result(20) => DANGLING_U35_Result_20,
       Result(21) => DANGLING_U35_Result_21,
       Result(22) => DANGLING_U35_Result_22,
       Result(23) => DANGLING_U35_Result_23,
       Result(24) => DANGLING_U35_Result_24,
       Result(25) => DANGLING_U35_Result_25,
       Result(26) => DANGLING_U35_Result_26,
       Result(27) => DANGLING_U35_Result_27,
       Result(28) => DANGLING_U35_Result_28,
       Result(29) => DANGLING_U35_Result_29,
       Result(30) => DANGLING_U35_Result_30,
       Result(31) => DANGLING_U35_Result_31,
       Result(32) => DANGLING_U35_Result_32,
       Result(33) => DANGLING_U35_Result_33,
       Result(34) => DANGLING_U35_Result_34,
       Result(35) => DANGLING_U35_Result_35,
       Result(36) => DANGLING_U35_Result_36,
       Result(37) => DANGLING_U35_Result_37,
       Result(38) => DANGLING_U35_Result_38,
       Result(39) => DANGLING_U35_Result_39,
       Result(40) => DANGLING_U35_Result_40,
       Result(41) => DANGLING_U35_Result_41,
       Result(42) => DANGLING_U35_Result_42,
       Result(43) => DANGLING_U35_Result_43,
       Result(44) => DANGLING_U35_Result_44,
       Result(45) => DANGLING_U35_Result_45,
       Result(46) => DANGLING_U35_Result_46,
       Result(47) => DANGLING_U35_Result_47,
       Result(48) => DANGLING_U35_Result_48,
       Result(49) => DANGLING_U35_Result_49,
       Result(50) => DANGLING_U35_Result_50,
       Result(51) => DANGLING_U35_Result_51,
       Result(52) => DANGLING_U35_Result_52,
       Result(53) => DANGLING_U35_Result_53,
       Result(54) => DANGLING_U35_Result_54,
       Result(55) => DANGLING_U35_Result_55,
       Result(56) => DANGLING_U35_Result_56,
       Result(57) => DANGLING_U35_Result_57,
       Result(58) => DANGLING_U35_Result_58,
       Result(59) => DANGLING_U35_Result_59,
       Result(60) => DANGLING_U35_Result_60,
       Result(61) => DANGLING_U35_Result_61,
       Result(62) => DANGLING_U35_Result_62,
       Result(63) => DANGLING_U35_Result_63,
       Result(64) => DANGLING_U35_Result_64,
       Result(65) => DANGLING_U35_Result_65,
       Result(66) => DANGLING_U35_Result_66,
       Result(67) => DANGLING_U35_Result_67,
       Result(68) => DANGLING_U35_Result_68,
       Result(69) => DANGLING_U35_Result_69,
       Result(70) => DANGLING_U35_Result_70,
       Result(71) => DANGLING_U35_Result_71,
       Result(72) => DANGLING_U35_Result_72,
       Result(73) => DANGLING_U35_Result_73,
       Result(74) => DANGLING_U35_Result_74,
       Result(75) => DANGLING_U35_Result_75,
       Result(76) => DANGLING_U35_Result_76,
       Result(77) => DANGLING_U35_Result_77,
       Result(78) => DANGLING_U35_Result_78,
       Result(79) => DANGLING_U35_Result_79,
       Result(80) => DANGLING_U35_Result_80,
       Result(81) => DANGLING_U35_Result_81,
       Result(82) => DANGLING_U35_Result_82,
       Result(83) => DANGLING_U35_Result_83,
       Result(84) => DANGLING_U35_Result_84,
       Result(85) => DANGLING_U35_Result_85,
       Result(86) => DANGLING_U35_Result_86,
       Result(87) => DANGLING_U35_Result_87,
       Result(88) => DANGLING_U35_Result_88,
       Result(89) => DANGLING_U35_Result_89,
       Result(90) => DANGLING_U35_Result_90,
       Result(91) => DANGLING_U35_Result_91,
       Result(92) => DANGLING_U35_Result_92,
       Result(93) => DANGLING_U35_Result_93,
       Result(94) => DANGLING_U35_Result_94,
       Result(95) => DANGLING_U35_Result_95,
       Result(96) => DANGLING_U35_Result_96,
       Result(97) => DANGLING_U35_Result_97,
       Result(98) => DANGLING_U35_Result_98,
       Result(99) => DANGLING_U35_Result_99,
       Result(100) => DANGLING_U35_Result_100,
       Result(101) => DANGLING_U35_Result_101,
       Result(102) => DANGLING_U35_Result_102,
       Result(103) => DANGLING_U35_Result_103,
       Result(104) => DANGLING_U35_Result_104,
       Result(105) => DANGLING_U35_Result_105,
       Result(106) => DANGLING_U35_Result_106,
       Result(107) => DANGLING_U35_Result_107,
       Result(108) => DANGLING_U35_Result_108,
       Result(109) => DANGLING_U35_Result_109,
       Result(110) => DANGLING_U35_Result_110,
       Result(111) => DANGLING_U35_Result_111,
       Result(112) => DANGLING_U35_Result_112,
       Result(113) => DANGLING_U35_Result_113,
       Result(114) => DANGLING_U35_Result_114,
       Result(115) => DANGLING_U35_Result_115,
       Result(116) => DANGLING_U35_Result_116,
       Result(117) => DANGLING_U35_Result_117,
       Result(118) => DANGLING_U35_Result_118,
       Result(119) => DANGLING_U35_Result_119,
       Result(120) => BUS2032(0),
       Result(121) => BUS2032(1),
       Result(122) => BUS2032(2),
       Result(123) => BUS2032(3),
       Result(124) => BUS2032(4),
       Result(125) => BUS2032(5),
       Result(126) => BUS2032(6),
       Result(127) => BUS2032(7),
       op_sel => BUS620
  );

U36 : byte_unit
  port map(
       A => BUS328,
       B => BUS297,
       Result => BUS209,
       op_sel => BUS616
  );

U37 : even_pipe_reg
  port map(
       Latency_d => BUS1961,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => NET600,
       RegdDst_d => BUS608,
       Unit_d(0) => BUS245(5),
       Unit_d(1) => BUS245(6),
       Unit_d(2) => BUS245(7),
       clk => Dangling_Input_Signal
  );

U39 : register_file
  port map(
       A_rd_addr => BUS1766,
       A_rd_data => BUS328,
       A_wr_addr => A_wr_addr,
       A_wr_data => A_wr_data,
       A_wr_en => A_wr_en,
       B_rd_addr => BUS1770,
       B_rd_data => BUS297,
       B_wr_addr => B_wr_addr,
       B_wr_data => B_wr_data,
       B_wr_en => B_wr_en,
       C_rd_addr => BUS1774,
       C_rd_data => BUS648,
       D_rd_addr => BUS1778,
       D_rd_data => BUS751,
       E_rd_addr => BUS1782,
       E_rd_data => BUS779,
       F_rd_addr(0) => BUS1786(1),
       F_rd_addr(1) => BUS1786(2),
       F_rd_addr(2) => BUS1786(3),
       F_rd_addr(3) => BUS1786(4),
       F_rd_addr(4) => BUS1786(5),
       F_rd_addr(5) => BUS1786(6),
       F_rd_addr(6) => BUS1786(7),
       F_rd_data => BUS789,
       clk => Dangling_Input_Signal
  );

U40 : permute_unit
  port map(
       A => BUS751,
       Result => BUS678,
       op_sel => BUS725
  );

U41 : branch_unit
  port map(
       A => BUS751,
       I16 => BUS772,
       PC => BUS741,
       Result => BUS686,
       T => BUS789,
       op_sel => BUS733
  );

U42 : local_store_unit
  port map(
       A => BUS751,
       B => BUS779,
       I10 => BUS762,
       I16 => BUS772,
       Result => BUS694,
       T => BUS789,
       clk => Dangling_Input_Signal,
       op_sel => BUS758
  );

U44 : odd_pipe_reg
  port map(
       Branch_d => NET1711,
       Latency_d => BUS1719,
       RegWr_d => NET1703,
       RegdDst_d => BUS1695,
       Result_d => BUS670,
       Unit_d => BUS709,
       clk => Dangling_Input_Signal
  );

U45 : even_pipe_reg
  port map(
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U46 : even_pipe_reg
  port map(
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U47 : even_pipe_reg
  port map(
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U48 : even_pipe_reg
  port map(
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U49 : even_pipe_reg
  port map(
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U50 : even_pipe_reg
  port map(
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U51 : odd_pipe_reg
  port map(
       Branch_d => Dangling_Input_Signal,
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U52 : odd_pipe_reg
  port map(
       Branch_d => Dangling_Input_Signal,
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U53 : odd_pipe_reg
  port map(
       Branch_d => Dangling_Input_Signal,
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U54 : odd_pipe_reg
  port map(
       Branch_d => Dangling_Input_Signal,
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U55 : odd_pipe_reg
  port map(
       Branch_d => Dangling_Input_Signal,
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U56 : odd_pipe_reg
  port map(
       Branch_d => Dangling_Input_Signal,
       Latency_d(0) => Dangling_Input_Signal,
       Latency_d(1) => Dangling_Input_Signal,
       Latency_d(2) => Dangling_Input_Signal,
       RegdDst_d(0) => Dangling_Input_Signal,
       RegdDst_d(1) => Dangling_Input_Signal,
       RegdDst_d(2) => Dangling_Input_Signal,
       RegdDst_d(3) => Dangling_Input_Signal,
       RegdDst_d(4) => Dangling_Input_Signal,
       RegdDst_d(5) => Dangling_Input_Signal,
       RegdDst_d(6) => Dangling_Input_Signal,
       Result_d(0) => Dangling_Input_Signal,
       Result_d(1) => Dangling_Input_Signal,
       Result_d(2) => Dangling_Input_Signal,
       Result_d(3) => Dangling_Input_Signal,
       Result_d(4) => Dangling_Input_Signal,
       Result_d(5) => Dangling_Input_Signal,
       Result_d(6) => Dangling_Input_Signal,
       Result_d(7) => Dangling_Input_Signal,
       Result_d(8) => Dangling_Input_Signal,
       Result_d(9) => Dangling_Input_Signal,
       Result_d(10) => Dangling_Input_Signal,
       Result_d(11) => Dangling_Input_Signal,
       Result_d(12) => Dangling_Input_Signal,
       Result_d(13) => Dangling_Input_Signal,
       Result_d(14) => Dangling_Input_Signal,
       Result_d(15) => Dangling_Input_Signal,
       Result_d(16) => Dangling_Input_Signal,
       Result_d(17) => Dangling_Input_Signal,
       Result_d(18) => Dangling_Input_Signal,
       Result_d(19) => Dangling_Input_Signal,
       Result_d(20) => Dangling_Input_Signal,
       Result_d(21) => Dangling_Input_Signal,
       Result_d(22) => Dangling_Input_Signal,
       Result_d(23) => Dangling_Input_Signal,
       Result_d(24) => Dangling_Input_Signal,
       Result_d(25) => Dangling_Input_Signal,
       Result_d(26) => Dangling_Input_Signal,
       Result_d(27) => Dangling_Input_Signal,
       Result_d(28) => Dangling_Input_Signal,
       Result_d(29) => Dangling_Input_Signal,
       Result_d(30) => Dangling_Input_Signal,
       Result_d(31) => Dangling_Input_Signal,
       Result_d(32) => Dangling_Input_Signal,
       Result_d(33) => Dangling_Input_Signal,
       Result_d(34) => Dangling_Input_Signal,
       Result_d(35) => Dangling_Input_Signal,
       Result_d(36) => Dangling_Input_Signal,
       Result_d(37) => Dangling_Input_Signal,
       Result_d(38) => Dangling_Input_Signal,
       Result_d(39) => Dangling_Input_Signal,
       Result_d(40) => Dangling_Input_Signal,
       Result_d(41) => Dangling_Input_Signal,
       Result_d(42) => Dangling_Input_Signal,
       Result_d(43) => Dangling_Input_Signal,
       Result_d(44) => Dangling_Input_Signal,
       Result_d(45) => Dangling_Input_Signal,
       Result_d(46) => Dangling_Input_Signal,
       Result_d(47) => Dangling_Input_Signal,
       Result_d(48) => Dangling_Input_Signal,
       Result_d(49) => Dangling_Input_Signal,
       Result_d(50) => Dangling_Input_Signal,
       Result_d(51) => Dangling_Input_Signal,
       Result_d(52) => Dangling_Input_Signal,
       Result_d(53) => Dangling_Input_Signal,
       Result_d(54) => Dangling_Input_Signal,
       Result_d(55) => Dangling_Input_Signal,
       Result_d(56) => Dangling_Input_Signal,
       Result_d(57) => Dangling_Input_Signal,
       Result_d(58) => Dangling_Input_Signal,
       Result_d(59) => Dangling_Input_Signal,
       Result_d(60) => Dangling_Input_Signal,
       Result_d(61) => Dangling_Input_Signal,
       Result_d(62) => Dangling_Input_Signal,
       Result_d(63) => Dangling_Input_Signal,
       Result_d(64) => Dangling_Input_Signal,
       Result_d(65) => Dangling_Input_Signal,
       Result_d(66) => Dangling_Input_Signal,
       Result_d(67) => Dangling_Input_Signal,
       Result_d(68) => Dangling_Input_Signal,
       Result_d(69) => Dangling_Input_Signal,
       Result_d(70) => Dangling_Input_Signal,
       Result_d(71) => Dangling_Input_Signal,
       Result_d(72) => Dangling_Input_Signal,
       Result_d(73) => Dangling_Input_Signal,
       Result_d(74) => Dangling_Input_Signal,
       Result_d(75) => Dangling_Input_Signal,
       Result_d(76) => Dangling_Input_Signal,
       Result_d(77) => Dangling_Input_Signal,
       Result_d(78) => Dangling_Input_Signal,
       Result_d(79) => Dangling_Input_Signal,
       Result_d(80) => Dangling_Input_Signal,
       Result_d(81) => Dangling_Input_Signal,
       Result_d(82) => Dangling_Input_Signal,
       Result_d(83) => Dangling_Input_Signal,
       Result_d(84) => Dangling_Input_Signal,
       Result_d(85) => Dangling_Input_Signal,
       Result_d(86) => Dangling_Input_Signal,
       Result_d(87) => Dangling_Input_Signal,
       Result_d(88) => Dangling_Input_Signal,
       Result_d(89) => Dangling_Input_Signal,
       Result_d(90) => Dangling_Input_Signal,
       Result_d(91) => Dangling_Input_Signal,
       Result_d(92) => Dangling_Input_Signal,
       Result_d(93) => Dangling_Input_Signal,
       Result_d(94) => Dangling_Input_Signal,
       Result_d(95) => Dangling_Input_Signal,
       Result_d(96) => Dangling_Input_Signal,
       Result_d(97) => Dangling_Input_Signal,
       Result_d(98) => Dangling_Input_Signal,
       Result_d(99) => Dangling_Input_Signal,
       Result_d(100) => Dangling_Input_Signal,
       Result_d(101) => Dangling_Input_Signal,
       Result_d(102) => Dangling_Input_Signal,
       Result_d(103) => Dangling_Input_Signal,
       Result_d(104) => Dangling_Input_Signal,
       Result_d(105) => Dangling_Input_Signal,
       Result_d(106) => Dangling_Input_Signal,
       Result_d(107) => Dangling_Input_Signal,
       Result_d(108) => Dangling_Input_Signal,
       Result_d(109) => Dangling_Input_Signal,
       Result_d(110) => Dangling_Input_Signal,
       Result_d(111) => Dangling_Input_Signal,
       Result_d(112) => Dangling_Input_Signal,
       Result_d(113) => Dangling_Input_Signal,
       Result_d(114) => Dangling_Input_Signal,
       Result_d(115) => Dangling_Input_Signal,
       Result_d(116) => Dangling_Input_Signal,
       Result_d(117) => Dangling_Input_Signal,
       Result_d(118) => Dangling_Input_Signal,
       Result_d(119) => Dangling_Input_Signal,
       Result_d(120) => Dangling_Input_Signal,
       Result_d(121) => Dangling_Input_Signal,
       Result_d(122) => Dangling_Input_Signal,
       Result_d(123) => Dangling_Input_Signal,
       Result_d(124) => Dangling_Input_Signal,
       Result_d(125) => Dangling_Input_Signal,
       Result_d(126) => Dangling_Input_Signal,
       Result_d(127) => Dangling_Input_Signal,
       RegWr_d => Dangling_Input_Signal,
       Unit_d(0) => Dangling_Input_Signal,
       Unit_d(1) => Dangling_Input_Signal,
       Unit_d(2) => Dangling_Input_Signal,
       clk => Dangling_Input_Signal
  );

U6 : forwarding_unit
  port map(
       A_reg(0) => Dangling_Input_Signal,
       A_reg(1) => Dangling_Input_Signal,
       A_reg(2) => Dangling_Input_Signal,
       A_reg(3) => Dangling_Input_Signal,
       A_reg(4) => Dangling_Input_Signal,
       A_reg(5) => Dangling_Input_Signal,
       A_reg(6) => Dangling_Input_Signal,
       A_reg(7) => Dangling_Input_Signal,
       A_reg(8) => Dangling_Input_Signal,
       A_reg(9) => Dangling_Input_Signal,
       A_reg(10) => Dangling_Input_Signal,
       A_reg(11) => Dangling_Input_Signal,
       A_reg(12) => Dangling_Input_Signal,
       A_reg(13) => Dangling_Input_Signal,
       A_reg(14) => Dangling_Input_Signal,
       A_reg(15) => Dangling_Input_Signal,
       A_reg(16) => Dangling_Input_Signal,
       A_reg(17) => Dangling_Input_Signal,
       A_reg(18) => Dangling_Input_Signal,
       A_reg(19) => Dangling_Input_Signal,
       A_reg(20) => Dangling_Input_Signal,
       A_reg(21) => Dangling_Input_Signal,
       A_reg(22) => Dangling_Input_Signal,
       A_reg(23) => Dangling_Input_Signal,
       A_reg(24) => Dangling_Input_Signal,
       A_reg(25) => Dangling_Input_Signal,
       A_reg(26) => Dangling_Input_Signal,
       A_reg(27) => Dangling_Input_Signal,
       A_reg(28) => Dangling_Input_Signal,
       A_reg(29) => Dangling_Input_Signal,
       A_reg(30) => Dangling_Input_Signal,
       A_reg(31) => Dangling_Input_Signal,
       A_reg(32) => Dangling_Input_Signal,
       A_reg(33) => Dangling_Input_Signal,
       A_reg(34) => Dangling_Input_Signal,
       A_reg(35) => Dangling_Input_Signal,
       A_reg(36) => Dangling_Input_Signal,
       A_reg(37) => Dangling_Input_Signal,
       A_reg(38) => Dangling_Input_Signal,
       A_reg(39) => Dangling_Input_Signal,
       A_reg(40) => Dangling_Input_Signal,
       A_reg(41) => Dangling_Input_Signal,
       A_reg(42) => Dangling_Input_Signal,
       A_reg(43) => Dangling_Input_Signal,
       A_reg(44) => Dangling_Input_Signal,
       A_reg(45) => Dangling_Input_Signal,
       A_reg(46) => Dangling_Input_Signal,
       A_reg(47) => Dangling_Input_Signal,
       A_reg(48) => Dangling_Input_Signal,
       A_reg(49) => Dangling_Input_Signal,
       A_reg(50) => Dangling_Input_Signal,
       A_reg(51) => Dangling_Input_Signal,
       A_reg(52) => Dangling_Input_Signal,
       A_reg(53) => Dangling_Input_Signal,
       A_reg(54) => Dangling_Input_Signal,
       A_reg(55) => Dangling_Input_Signal,
       A_reg(56) => Dangling_Input_Signal,
       A_reg(57) => Dangling_Input_Signal,
       A_reg(58) => Dangling_Input_Signal,
       A_reg(59) => Dangling_Input_Signal,
       A_reg(60) => Dangling_Input_Signal,
       A_reg(61) => Dangling_Input_Signal,
       A_reg(62) => Dangling_Input_Signal,
       A_reg(63) => Dangling_Input_Signal,
       A_reg(64) => Dangling_Input_Signal,
       A_reg(65) => Dangling_Input_Signal,
       A_reg(66) => Dangling_Input_Signal,
       A_reg(67) => Dangling_Input_Signal,
       A_reg(68) => Dangling_Input_Signal,
       A_reg(69) => Dangling_Input_Signal,
       A_reg(70) => Dangling_Input_Signal,
       A_reg(71) => Dangling_Input_Signal,
       A_reg(72) => Dangling_Input_Signal,
       A_reg(73) => Dangling_Input_Signal,
       A_reg(74) => Dangling_Input_Signal,
       A_reg(75) => Dangling_Input_Signal,
       A_reg(76) => Dangling_Input_Signal,
       A_reg(77) => Dangling_Input_Signal,
       A_reg(78) => Dangling_Input_Signal,
       A_reg(79) => Dangling_Input_Signal,
       A_reg(80) => Dangling_Input_Signal,
       A_reg(81) => Dangling_Input_Signal,
       A_reg(82) => Dangling_Input_Signal,
       A_reg(83) => Dangling_Input_Signal,
       A_reg(84) => Dangling_Input_Signal,
       A_reg(85) => Dangling_Input_Signal,
       A_reg(86) => Dangling_Input_Signal,
       A_reg(87) => Dangling_Input_Signal,
       A_reg(88) => Dangling_Input_Signal,
       A_reg(89) => Dangling_Input_Signal,
       A_reg(90) => Dangling_Input_Signal,
       A_reg(91) => Dangling_Input_Signal,
       A_reg(92) => Dangling_Input_Signal,
       A_reg(93) => Dangling_Input_Signal,
       A_reg(94) => Dangling_Input_Signal,
       A_reg(95) => Dangling_Input_Signal,
       A_reg(96) => Dangling_Input_Signal,
       A_reg(97) => Dangling_Input_Signal,
       A_reg(98) => Dangling_Input_Signal,
       A_reg(99) => Dangling_Input_Signal,
       A_reg(100) => Dangling_Input_Signal,
       A_reg(101) => Dangling_Input_Signal,
       A_reg(102) => Dangling_Input_Signal,
       A_reg(103) => Dangling_Input_Signal,
       A_reg(104) => Dangling_Input_Signal,
       A_reg(105) => Dangling_Input_Signal,
       A_reg(106) => Dangling_Input_Signal,
       A_reg(107) => Dangling_Input_Signal,
       A_reg(108) => Dangling_Input_Signal,
       A_reg(109) => Dangling_Input_Signal,
       A_reg(110) => Dangling_Input_Signal,
       A_reg(111) => Dangling_Input_Signal,
       A_reg(112) => Dangling_Input_Signal,
       A_reg(113) => Dangling_Input_Signal,
       A_reg(114) => Dangling_Input_Signal,
       A_reg(115) => Dangling_Input_Signal,
       A_reg(116) => Dangling_Input_Signal,
       A_reg(117) => Dangling_Input_Signal,
       A_reg(118) => Dangling_Input_Signal,
       A_reg(119) => Dangling_Input_Signal,
       A_reg(120) => Dangling_Input_Signal,
       A_reg(121) => Dangling_Input_Signal,
       A_reg(122) => Dangling_Input_Signal,
       A_reg(123) => Dangling_Input_Signal,
       A_reg(124) => Dangling_Input_Signal,
       A_reg(125) => Dangling_Input_Signal,
       A_reg(126) => Dangling_Input_Signal,
       A_reg(127) => Dangling_Input_Signal,
       B_reg(0) => Dangling_Input_Signal,
       B_reg(1) => Dangling_Input_Signal,
       B_reg(2) => Dangling_Input_Signal,
       B_reg(3) => Dangling_Input_Signal,
       B_reg(4) => Dangling_Input_Signal,
       B_reg(5) => Dangling_Input_Signal,
       B_reg(6) => Dangling_Input_Signal,
       B_reg(7) => Dangling_Input_Signal,
       B_reg(8) => Dangling_Input_Signal,
       B_reg(9) => Dangling_Input_Signal,
       B_reg(10) => Dangling_Input_Signal,
       B_reg(11) => Dangling_Input_Signal,
       B_reg(12) => Dangling_Input_Signal,
       B_reg(13) => Dangling_Input_Signal,
       B_reg(14) => Dangling_Input_Signal,
       B_reg(15) => Dangling_Input_Signal,
       B_reg(16) => Dangling_Input_Signal,
       B_reg(17) => Dangling_Input_Signal,
       B_reg(18) => Dangling_Input_Signal,
       B_reg(19) => Dangling_Input_Signal,
       B_reg(20) => Dangling_Input_Signal,
       B_reg(21) => Dangling_Input_Signal,
       B_reg(22) => Dangling_Input_Signal,
       B_reg(23) => Dangling_Input_Signal,
       B_reg(24) => Dangling_Input_Signal,
       B_reg(25) => Dangling_Input_Signal,
       B_reg(26) => Dangling_Input_Signal,
       B_reg(27) => Dangling_Input_Signal,
       B_reg(28) => Dangling_Input_Signal,
       B_reg(29) => Dangling_Input_Signal,
       B_reg(30) => Dangling_Input_Signal,
       B_reg(31) => Dangling_Input_Signal,
       B_reg(32) => Dangling_Input_Signal,
       B_reg(33) => Dangling_Input_Signal,
       B_reg(34) => Dangling_Input_Signal,
       B_reg(35) => Dangling_Input_Signal,
       B_reg(36) => Dangling_Input_Signal,
       B_reg(37) => Dangling_Input_Signal,
       B_reg(38) => Dangling_Input_Signal,
       B_reg(39) => Dangling_Input_Signal,
       B_reg(40) => Dangling_Input_Signal,
       B_reg(41) => Dangling_Input_Signal,
       B_reg(42) => Dangling_Input_Signal,
       B_reg(43) => Dangling_Input_Signal,
       B_reg(44) => Dangling_Input_Signal,
       B_reg(45) => Dangling_Input_Signal,
       B_reg(46) => Dangling_Input_Signal,
       B_reg(47) => Dangling_Input_Signal,
       B_reg(48) => Dangling_Input_Signal,
       B_reg(49) => Dangling_Input_Signal,
       B_reg(50) => Dangling_Input_Signal,
       B_reg(51) => Dangling_Input_Signal,
       B_reg(52) => Dangling_Input_Signal,
       B_reg(53) => Dangling_Input_Signal,
       B_reg(54) => Dangling_Input_Signal,
       B_reg(55) => Dangling_Input_Signal,
       B_reg(56) => Dangling_Input_Signal,
       B_reg(57) => Dangling_Input_Signal,
       B_reg(58) => Dangling_Input_Signal,
       B_reg(59) => Dangling_Input_Signal,
       B_reg(60) => Dangling_Input_Signal,
       B_reg(61) => Dangling_Input_Signal,
       B_reg(62) => Dangling_Input_Signal,
       B_reg(63) => Dangling_Input_Signal,
       B_reg(64) => Dangling_Input_Signal,
       B_reg(65) => Dangling_Input_Signal,
       B_reg(66) => Dangling_Input_Signal,
       B_reg(67) => Dangling_Input_Signal,
       B_reg(68) => Dangling_Input_Signal,
       B_reg(69) => Dangling_Input_Signal,
       B_reg(70) => Dangling_Input_Signal,
       B_reg(71) => Dangling_Input_Signal,
       B_reg(72) => Dangling_Input_Signal,
       B_reg(73) => Dangling_Input_Signal,
       B_reg(74) => Dangling_Input_Signal,
       B_reg(75) => Dangling_Input_Signal,
       B_reg(76) => Dangling_Input_Signal,
       B_reg(77) => Dangling_Input_Signal,
       B_reg(78) => Dangling_Input_Signal,
       B_reg(79) => Dangling_Input_Signal,
       B_reg(80) => Dangling_Input_Signal,
       B_reg(81) => Dangling_Input_Signal,
       B_reg(82) => Dangling_Input_Signal,
       B_reg(83) => Dangling_Input_Signal,
       B_reg(84) => Dangling_Input_Signal,
       B_reg(85) => Dangling_Input_Signal,
       B_reg(86) => Dangling_Input_Signal,
       B_reg(87) => Dangling_Input_Signal,
       B_reg(88) => Dangling_Input_Signal,
       B_reg(89) => Dangling_Input_Signal,
       B_reg(90) => Dangling_Input_Signal,
       B_reg(91) => Dangling_Input_Signal,
       B_reg(92) => Dangling_Input_Signal,
       B_reg(93) => Dangling_Input_Signal,
       B_reg(94) => Dangling_Input_Signal,
       B_reg(95) => Dangling_Input_Signal,
       B_reg(96) => Dangling_Input_Signal,
       B_reg(97) => Dangling_Input_Signal,
       B_reg(98) => Dangling_Input_Signal,
       B_reg(99) => Dangling_Input_Signal,
       B_reg(100) => Dangling_Input_Signal,
       B_reg(101) => Dangling_Input_Signal,
       B_reg(102) => Dangling_Input_Signal,
       B_reg(103) => Dangling_Input_Signal,
       B_reg(104) => Dangling_Input_Signal,
       B_reg(105) => Dangling_Input_Signal,
       B_reg(106) => Dangling_Input_Signal,
       B_reg(107) => Dangling_Input_Signal,
       B_reg(108) => Dangling_Input_Signal,
       B_reg(109) => Dangling_Input_Signal,
       B_reg(110) => Dangling_Input_Signal,
       B_reg(111) => Dangling_Input_Signal,
       B_reg(112) => Dangling_Input_Signal,
       B_reg(113) => Dangling_Input_Signal,
       B_reg(114) => Dangling_Input_Signal,
       B_reg(115) => Dangling_Input_Signal,
       B_reg(116) => Dangling_Input_Signal,
       B_reg(117) => Dangling_Input_Signal,
       B_reg(118) => Dangling_Input_Signal,
       B_reg(119) => Dangling_Input_Signal,
       B_reg(120) => Dangling_Input_Signal,
       B_reg(121) => Dangling_Input_Signal,
       B_reg(122) => Dangling_Input_Signal,
       B_reg(123) => Dangling_Input_Signal,
       B_reg(124) => Dangling_Input_Signal,
       B_reg(125) => Dangling_Input_Signal,
       B_reg(126) => Dangling_Input_Signal,
       B_reg(127) => Dangling_Input_Signal,
       C_reg(0) => Dangling_Input_Signal,
       C_reg(1) => Dangling_Input_Signal,
       C_reg(2) => Dangling_Input_Signal,
       C_reg(3) => Dangling_Input_Signal,
       C_reg(4) => Dangling_Input_Signal,
       C_reg(5) => Dangling_Input_Signal,
       C_reg(6) => Dangling_Input_Signal,
       C_reg(7) => Dangling_Input_Signal,
       C_reg(8) => Dangling_Input_Signal,
       C_reg(9) => Dangling_Input_Signal,
       C_reg(10) => Dangling_Input_Signal,
       C_reg(11) => Dangling_Input_Signal,
       C_reg(12) => Dangling_Input_Signal,
       C_reg(13) => Dangling_Input_Signal,
       C_reg(14) => Dangling_Input_Signal,
       C_reg(15) => Dangling_Input_Signal,
       C_reg(16) => Dangling_Input_Signal,
       C_reg(17) => Dangling_Input_Signal,
       C_reg(18) => Dangling_Input_Signal,
       C_reg(19) => Dangling_Input_Signal,
       C_reg(20) => Dangling_Input_Signal,
       C_reg(21) => Dangling_Input_Signal,
       C_reg(22) => Dangling_Input_Signal,
       C_reg(23) => Dangling_Input_Signal,
       C_reg(24) => Dangling_Input_Signal,
       C_reg(25) => Dangling_Input_Signal,
       C_reg(26) => Dangling_Input_Signal,
       C_reg(27) => Dangling_Input_Signal,
       C_reg(28) => Dangling_Input_Signal,
       C_reg(29) => Dangling_Input_Signal,
       C_reg(30) => Dangling_Input_Signal,
       C_reg(31) => Dangling_Input_Signal,
       C_reg(32) => Dangling_Input_Signal,
       C_reg(33) => Dangling_Input_Signal,
       C_reg(34) => Dangling_Input_Signal,
       C_reg(35) => Dangling_Input_Signal,
       C_reg(36) => Dangling_Input_Signal,
       C_reg(37) => Dangling_Input_Signal,
       C_reg(38) => Dangling_Input_Signal,
       C_reg(39) => Dangling_Input_Signal,
       C_reg(40) => Dangling_Input_Signal,
       C_reg(41) => Dangling_Input_Signal,
       C_reg(42) => Dangling_Input_Signal,
       C_reg(43) => Dangling_Input_Signal,
       C_reg(44) => Dangling_Input_Signal,
       C_reg(45) => Dangling_Input_Signal,
       C_reg(46) => Dangling_Input_Signal,
       C_reg(47) => Dangling_Input_Signal,
       C_reg(48) => Dangling_Input_Signal,
       C_reg(49) => Dangling_Input_Signal,
       C_reg(50) => Dangling_Input_Signal,
       C_reg(51) => Dangling_Input_Signal,
       C_reg(52) => Dangling_Input_Signal,
       C_reg(53) => Dangling_Input_Signal,
       C_reg(54) => Dangling_Input_Signal,
       C_reg(55) => Dangling_Input_Signal,
       C_reg(56) => Dangling_Input_Signal,
       C_reg(57) => Dangling_Input_Signal,
       C_reg(58) => Dangling_Input_Signal,
       C_reg(59) => Dangling_Input_Signal,
       C_reg(60) => Dangling_Input_Signal,
       C_reg(61) => Dangling_Input_Signal,
       C_reg(62) => Dangling_Input_Signal,
       C_reg(63) => Dangling_Input_Signal,
       C_reg(64) => Dangling_Input_Signal,
       C_reg(65) => Dangling_Input_Signal,
       C_reg(66) => Dangling_Input_Signal,
       C_reg(67) => Dangling_Input_Signal,
       C_reg(68) => Dangling_Input_Signal,
       C_reg(69) => Dangling_Input_Signal,
       C_reg(70) => Dangling_Input_Signal,
       C_reg(71) => Dangling_Input_Signal,
       C_reg(72) => Dangling_Input_Signal,
       C_reg(73) => Dangling_Input_Signal,
       C_reg(74) => Dangling_Input_Signal,
       C_reg(75) => Dangling_Input_Signal,
       C_reg(76) => Dangling_Input_Signal,
       C_reg(77) => Dangling_Input_Signal,
       C_reg(78) => Dangling_Input_Signal,
       C_reg(79) => Dangling_Input_Signal,
       C_reg(80) => Dangling_Input_Signal,
       C_reg(81) => Dangling_Input_Signal,
       C_reg(82) => Dangling_Input_Signal,
       C_reg(83) => Dangling_Input_Signal,
       C_reg(84) => Dangling_Input_Signal,
       C_reg(85) => Dangling_Input_Signal,
       C_reg(86) => Dangling_Input_Signal,
       C_reg(87) => Dangling_Input_Signal,
       C_reg(88) => Dangling_Input_Signal,
       C_reg(89) => Dangling_Input_Signal,
       C_reg(90) => Dangling_Input_Signal,
       C_reg(91) => Dangling_Input_Signal,
       C_reg(92) => Dangling_Input_Signal,
       C_reg(93) => Dangling_Input_Signal,
       C_reg(94) => Dangling_Input_Signal,
       C_reg(95) => Dangling_Input_Signal,
       C_reg(96) => Dangling_Input_Signal,
       C_reg(97) => Dangling_Input_Signal,
       C_reg(98) => Dangling_Input_Signal,
       C_reg(99) => Dangling_Input_Signal,
       C_reg(100) => Dangling_Input_Signal,
       C_reg(101) => Dangling_Input_Signal,
       C_reg(102) => Dangling_Input_Signal,
       C_reg(103) => Dangling_Input_Signal,
       C_reg(104) => Dangling_Input_Signal,
       C_reg(105) => Dangling_Input_Signal,
       C_reg(106) => Dangling_Input_Signal,
       C_reg(107) => Dangling_Input_Signal,
       C_reg(108) => Dangling_Input_Signal,
       C_reg(109) => Dangling_Input_Signal,
       C_reg(110) => Dangling_Input_Signal,
       C_reg(111) => Dangling_Input_Signal,
       C_reg(112) => Dangling_Input_Signal,
       C_reg(113) => Dangling_Input_Signal,
       C_reg(114) => Dangling_Input_Signal,
       C_reg(115) => Dangling_Input_Signal,
       C_reg(116) => Dangling_Input_Signal,
       C_reg(117) => Dangling_Input_Signal,
       C_reg(118) => Dangling_Input_Signal,
       C_reg(119) => Dangling_Input_Signal,
       C_reg(120) => Dangling_Input_Signal,
       C_reg(121) => Dangling_Input_Signal,
       C_reg(122) => Dangling_Input_Signal,
       C_reg(123) => Dangling_Input_Signal,
       C_reg(124) => Dangling_Input_Signal,
       C_reg(125) => Dangling_Input_Signal,
       C_reg(126) => Dangling_Input_Signal,
       C_reg(127) => Dangling_Input_Signal,
       D_reg(0) => Dangling_Input_Signal,
       D_reg(1) => Dangling_Input_Signal,
       D_reg(2) => Dangling_Input_Signal,
       D_reg(3) => Dangling_Input_Signal,
       D_reg(4) => Dangling_Input_Signal,
       D_reg(5) => Dangling_Input_Signal,
       D_reg(6) => Dangling_Input_Signal,
       D_reg(7) => Dangling_Input_Signal,
       D_reg(8) => Dangling_Input_Signal,
       D_reg(9) => Dangling_Input_Signal,
       D_reg(10) => Dangling_Input_Signal,
       D_reg(11) => Dangling_Input_Signal,
       D_reg(12) => Dangling_Input_Signal,
       D_reg(13) => Dangling_Input_Signal,
       D_reg(14) => Dangling_Input_Signal,
       D_reg(15) => Dangling_Input_Signal,
       D_reg(16) => Dangling_Input_Signal,
       D_reg(17) => Dangling_Input_Signal,
       D_reg(18) => Dangling_Input_Signal,
       D_reg(19) => Dangling_Input_Signal,
       D_reg(20) => Dangling_Input_Signal,
       D_reg(21) => Dangling_Input_Signal,
       D_reg(22) => Dangling_Input_Signal,
       D_reg(23) => Dangling_Input_Signal,
       D_reg(24) => Dangling_Input_Signal,
       D_reg(25) => Dangling_Input_Signal,
       D_reg(26) => Dangling_Input_Signal,
       D_reg(27) => Dangling_Input_Signal,
       D_reg(28) => Dangling_Input_Signal,
       D_reg(29) => Dangling_Input_Signal,
       D_reg(30) => Dangling_Input_Signal,
       D_reg(31) => Dangling_Input_Signal,
       D_reg(32) => Dangling_Input_Signal,
       D_reg(33) => Dangling_Input_Signal,
       D_reg(34) => Dangling_Input_Signal,
       D_reg(35) => Dangling_Input_Signal,
       D_reg(36) => Dangling_Input_Signal,
       D_reg(37) => Dangling_Input_Signal,
       D_reg(38) => Dangling_Input_Signal,
       D_reg(39) => Dangling_Input_Signal,
       D_reg(40) => Dangling_Input_Signal,
       D_reg(41) => Dangling_Input_Signal,
       D_reg(42) => Dangling_Input_Signal,
       D_reg(43) => Dangling_Input_Signal,
       D_reg(44) => Dangling_Input_Signal,
       D_reg(45) => Dangling_Input_Signal,
       D_reg(46) => Dangling_Input_Signal,
       D_reg(47) => Dangling_Input_Signal,
       D_reg(48) => Dangling_Input_Signal,
       D_reg(49) => Dangling_Input_Signal,
       D_reg(50) => Dangling_Input_Signal,
       D_reg(51) => Dangling_Input_Signal,
       D_reg(52) => Dangling_Input_Signal,
       D_reg(53) => Dangling_Input_Signal,
       D_reg(54) => Dangling_Input_Signal,
       D_reg(55) => Dangling_Input_Signal,
       D_reg(56) => Dangling_Input_Signal,
       D_reg(57) => Dangling_Input_Signal,
       D_reg(58) => Dangling_Input_Signal,
       D_reg(59) => Dangling_Input_Signal,
       D_reg(60) => Dangling_Input_Signal,
       D_reg(61) => Dangling_Input_Signal,
       D_reg(62) => Dangling_Input_Signal,
       D_reg(63) => Dangling_Input_Signal,
       D_reg(64) => Dangling_Input_Signal,
       D_reg(65) => Dangling_Input_Signal,
       D_reg(66) => Dangling_Input_Signal,
       D_reg(67) => Dangling_Input_Signal,
       D_reg(68) => Dangling_Input_Signal,
       D_reg(69) => Dangling_Input_Signal,
       D_reg(70) => Dangling_Input_Signal,
       D_reg(71) => Dangling_Input_Signal,
       D_reg(72) => Dangling_Input_Signal,
       D_reg(73) => Dangling_Input_Signal,
       D_reg(74) => Dangling_Input_Signal,
       D_reg(75) => Dangling_Input_Signal,
       D_reg(76) => Dangling_Input_Signal,
       D_reg(77) => Dangling_Input_Signal,
       D_reg(78) => Dangling_Input_Signal,
       D_reg(79) => Dangling_Input_Signal,
       D_reg(80) => Dangling_Input_Signal,
       D_reg(81) => Dangling_Input_Signal,
       D_reg(82) => Dangling_Input_Signal,
       D_reg(83) => Dangling_Input_Signal,
       D_reg(84) => Dangling_Input_Signal,
       D_reg(85) => Dangling_Input_Signal,
       D_reg(86) => Dangling_Input_Signal,
       D_reg(87) => Dangling_Input_Signal,
       D_reg(88) => Dangling_Input_Signal,
       D_reg(89) => Dangling_Input_Signal,
       D_reg(90) => Dangling_Input_Signal,
       D_reg(91) => Dangling_Input_Signal,
       D_reg(92) => Dangling_Input_Signal,
       D_reg(93) => Dangling_Input_Signal,
       D_reg(94) => Dangling_Input_Signal,
       D_reg(95) => Dangling_Input_Signal,
       D_reg(96) => Dangling_Input_Signal,
       D_reg(97) => Dangling_Input_Signal,
       D_reg(98) => Dangling_Input_Signal,
       D_reg(99) => Dangling_Input_Signal,
       D_reg(100) => Dangling_Input_Signal,
       D_reg(101) => Dangling_Input_Signal,
       D_reg(102) => Dangling_Input_Signal,
       D_reg(103) => Dangling_Input_Signal,
       D_reg(104) => Dangling_Input_Signal,
       D_reg(105) => Dangling_Input_Signal,
       D_reg(106) => Dangling_Input_Signal,
       D_reg(107) => Dangling_Input_Signal,
       D_reg(108) => Dangling_Input_Signal,
       D_reg(109) => Dangling_Input_Signal,
       D_reg(110) => Dangling_Input_Signal,
       D_reg(111) => Dangling_Input_Signal,
       D_reg(112) => Dangling_Input_Signal,
       D_reg(113) => Dangling_Input_Signal,
       D_reg(114) => Dangling_Input_Signal,
       D_reg(115) => Dangling_Input_Signal,
       D_reg(116) => Dangling_Input_Signal,
       D_reg(117) => Dangling_Input_Signal,
       D_reg(118) => Dangling_Input_Signal,
       D_reg(119) => Dangling_Input_Signal,
       D_reg(120) => Dangling_Input_Signal,
       D_reg(121) => Dangling_Input_Signal,
       D_reg(122) => Dangling_Input_Signal,
       D_reg(123) => Dangling_Input_Signal,
       D_reg(124) => Dangling_Input_Signal,
       D_reg(125) => Dangling_Input_Signal,
       D_reg(126) => Dangling_Input_Signal,
       D_reg(127) => Dangling_Input_Signal,
       even1_Latency(0) => Dangling_Input_Signal,
       even1_Latency(1) => Dangling_Input_Signal,
       even1_Latency(2) => Dangling_Input_Signal,
       even1_RegDst(0) => Dangling_Input_Signal,
       even1_RegDst(1) => Dangling_Input_Signal,
       even1_RegDst(2) => Dangling_Input_Signal,
       even1_RegDst(3) => Dangling_Input_Signal,
       even1_RegDst(4) => Dangling_Input_Signal,
       even1_RegDst(5) => Dangling_Input_Signal,
       even1_RegDst(6) => Dangling_Input_Signal,
       even1_Result(0) => Dangling_Input_Signal,
       even1_Result(1) => Dangling_Input_Signal,
       even1_Result(2) => Dangling_Input_Signal,
       even1_Result(3) => Dangling_Input_Signal,
       even1_Result(4) => Dangling_Input_Signal,
       even1_Result(5) => Dangling_Input_Signal,
       even1_Result(6) => Dangling_Input_Signal,
       even1_Result(7) => Dangling_Input_Signal,
       even1_Result(8) => Dangling_Input_Signal,
       even1_Result(9) => Dangling_Input_Signal,
       even1_Result(10) => Dangling_Input_Signal,
       even1_Result(11) => Dangling_Input_Signal,
       even1_Result(12) => Dangling_Input_Signal,
       even1_Result(13) => Dangling_Input_Signal,
       even1_Result(14) => Dangling_Input_Signal,
       even1_Result(15) => Dangling_Input_Signal,
       even1_Result(16) => Dangling_Input_Signal,
       even1_Result(17) => Dangling_Input_Signal,
       even1_Result(18) => Dangling_Input_Signal,
       even1_Result(19) => Dangling_Input_Signal,
       even1_Result(20) => Dangling_Input_Signal,
       even1_Result(21) => Dangling_Input_Signal,
       even1_Result(22) => Dangling_Input_Signal,
       even1_Result(23) => Dangling_Input_Signal,
       even1_Result(24) => Dangling_Input_Signal,
       even1_Result(25) => Dangling_Input_Signal,
       even1_Result(26) => Dangling_Input_Signal,
       even1_Result(27) => Dangling_Input_Signal,
       even1_Result(28) => Dangling_Input_Signal,
       even1_Result(29) => Dangling_Input_Signal,
       even1_Result(30) => Dangling_Input_Signal,
       even1_Result(31) => Dangling_Input_Signal,
       even1_Result(32) => Dangling_Input_Signal,
       even1_Result(33) => Dangling_Input_Signal,
       even1_Result(34) => Dangling_Input_Signal,
       even1_Result(35) => Dangling_Input_Signal,
       even1_Result(36) => Dangling_Input_Signal,
       even1_Result(37) => Dangling_Input_Signal,
       even1_Result(38) => Dangling_Input_Signal,
       even1_Result(39) => Dangling_Input_Signal,
       even1_Result(40) => Dangling_Input_Signal,
       even1_Result(41) => Dangling_Input_Signal,
       even1_Result(42) => Dangling_Input_Signal,
       even1_Result(43) => Dangling_Input_Signal,
       even1_Result(44) => Dangling_Input_Signal,
       even1_Result(45) => Dangling_Input_Signal,
       even1_Result(46) => Dangling_Input_Signal,
       even1_Result(47) => Dangling_Input_Signal,
       even1_Result(48) => Dangling_Input_Signal,
       even1_Result(49) => Dangling_Input_Signal,
       even1_Result(50) => Dangling_Input_Signal,
       even1_Result(51) => Dangling_Input_Signal,
       even1_Result(52) => Dangling_Input_Signal,
       even1_Result(53) => Dangling_Input_Signal,
       even1_Result(54) => Dangling_Input_Signal,
       even1_Result(55) => Dangling_Input_Signal,
       even1_Result(56) => Dangling_Input_Signal,
       even1_Result(57) => Dangling_Input_Signal,
       even1_Result(58) => Dangling_Input_Signal,
       even1_Result(59) => Dangling_Input_Signal,
       even1_Result(60) => Dangling_Input_Signal,
       even1_Result(61) => Dangling_Input_Signal,
       even1_Result(62) => Dangling_Input_Signal,
       even1_Result(63) => Dangling_Input_Signal,
       even1_Result(64) => Dangling_Input_Signal,
       even1_Result(65) => Dangling_Input_Signal,
       even1_Result(66) => Dangling_Input_Signal,
       even1_Result(67) => Dangling_Input_Signal,
       even1_Result(68) => Dangling_Input_Signal,
       even1_Result(69) => Dangling_Input_Signal,
       even1_Result(70) => Dangling_Input_Signal,
       even1_Result(71) => Dangling_Input_Signal,
       even1_Result(72) => Dangling_Input_Signal,
       even1_Result(73) => Dangling_Input_Signal,
       even1_Result(74) => Dangling_Input_Signal,
       even1_Result(75) => Dangling_Input_Signal,
       even1_Result(76) => Dangling_Input_Signal,
       even1_Result(77) => Dangling_Input_Signal,
       even1_Result(78) => Dangling_Input_Signal,
       even1_Result(79) => Dangling_Input_Signal,
       even1_Result(80) => Dangling_Input_Signal,
       even1_Result(81) => Dangling_Input_Signal,
       even1_Result(82) => Dangling_Input_Signal,
       even1_Result(83) => Dangling_Input_Signal,
       even1_Result(84) => Dangling_Input_Signal,
       even1_Result(85) => Dangling_Input_Signal,
       even1_Result(86) => Dangling_Input_Signal,
       even1_Result(87) => Dangling_Input_Signal,
       even1_Result(88) => Dangling_Input_Signal,
       even1_Result(89) => Dangling_Input_Signal,
       even1_Result(90) => Dangling_Input_Signal,
       even1_Result(91) => Dangling_Input_Signal,
       even1_Result(92) => Dangling_Input_Signal,
       even1_Result(93) => Dangling_Input_Signal,
       even1_Result(94) => Dangling_Input_Signal,
       even1_Result(95) => Dangling_Input_Signal,
       even1_Result(96) => Dangling_Input_Signal,
       even1_Result(97) => Dangling_Input_Signal,
       even1_Result(98) => Dangling_Input_Signal,
       even1_Result(99) => Dangling_Input_Signal,
       even1_Result(100) => Dangling_Input_Signal,
       even1_Result(101) => Dangling_Input_Signal,
       even1_Result(102) => Dangling_Input_Signal,
       even1_Result(103) => Dangling_Input_Signal,
       even1_Result(104) => Dangling_Input_Signal,
       even1_Result(105) => Dangling_Input_Signal,
       even1_Result(106) => Dangling_Input_Signal,
       even1_Result(107) => Dangling_Input_Signal,
       even1_Result(108) => Dangling_Input_Signal,
       even1_Result(109) => Dangling_Input_Signal,
       even1_Result(110) => Dangling_Input_Signal,
       even1_Result(111) => Dangling_Input_Signal,
       even1_Result(112) => Dangling_Input_Signal,
       even1_Result(113) => Dangling_Input_Signal,
       even1_Result(114) => Dangling_Input_Signal,
       even1_Result(115) => Dangling_Input_Signal,
       even1_Result(116) => Dangling_Input_Signal,
       even1_Result(117) => Dangling_Input_Signal,
       even1_Result(118) => Dangling_Input_Signal,
       even1_Result(119) => Dangling_Input_Signal,
       even1_Result(120) => Dangling_Input_Signal,
       even1_Result(121) => Dangling_Input_Signal,
       even1_Result(122) => Dangling_Input_Signal,
       even1_Result(123) => Dangling_Input_Signal,
       even1_Result(124) => Dangling_Input_Signal,
       even1_Result(125) => Dangling_Input_Signal,
       even1_Result(126) => Dangling_Input_Signal,
       even1_Result(127) => Dangling_Input_Signal,
       even2_Latency(0) => Dangling_Input_Signal,
       even2_Latency(1) => Dangling_Input_Signal,
       even2_Latency(2) => Dangling_Input_Signal,
       even2_RegDst(0) => Dangling_Input_Signal,
       even2_RegDst(1) => Dangling_Input_Signal,
       even2_RegDst(2) => Dangling_Input_Signal,
       even2_RegDst(3) => Dangling_Input_Signal,
       even2_RegDst(4) => Dangling_Input_Signal,
       even2_RegDst(5) => Dangling_Input_Signal,
       even2_RegDst(6) => Dangling_Input_Signal,
       even2_Result(0) => Dangling_Input_Signal,
       even2_Result(1) => Dangling_Input_Signal,
       even2_Result(2) => Dangling_Input_Signal,
       even2_Result(3) => Dangling_Input_Signal,
       even2_Result(4) => Dangling_Input_Signal,
       even2_Result(5) => Dangling_Input_Signal,
       even2_Result(6) => Dangling_Input_Signal,
       even2_Result(7) => Dangling_Input_Signal,
       even2_Result(8) => Dangling_Input_Signal,
       even2_Result(9) => Dangling_Input_Signal,
       even2_Result(10) => Dangling_Input_Signal,
       even2_Result(11) => Dangling_Input_Signal,
       even2_Result(12) => Dangling_Input_Signal,
       even2_Result(13) => Dangling_Input_Signal,
       even2_Result(14) => Dangling_Input_Signal,
       even2_Result(15) => Dangling_Input_Signal,
       even2_Result(16) => Dangling_Input_Signal,
       even2_Result(17) => Dangling_Input_Signal,
       even2_Result(18) => Dangling_Input_Signal,
       even2_Result(19) => Dangling_Input_Signal,
       even2_Result(20) => Dangling_Input_Signal,
       even2_Result(21) => Dangling_Input_Signal,
       even2_Result(22) => Dangling_Input_Signal,
       even2_Result(23) => Dangling_Input_Signal,
       even2_Result(24) => Dangling_Input_Signal,
       even2_Result(25) => Dangling_Input_Signal,
       even2_Result(26) => Dangling_Input_Signal,
       even2_Result(27) => Dangling_Input_Signal,
       even2_Result(28) => Dangling_Input_Signal,
       even2_Result(29) => Dangling_Input_Signal,
       even2_Result(30) => Dangling_Input_Signal,
       even2_Result(31) => Dangling_Input_Signal,
       even2_Result(32) => Dangling_Input_Signal,
       even2_Result(33) => Dangling_Input_Signal,
       even2_Result(34) => Dangling_Input_Signal,
       even2_Result(35) => Dangling_Input_Signal,
       even2_Result(36) => Dangling_Input_Signal,
       even2_Result(37) => Dangling_Input_Signal,
       even2_Result(38) => Dangling_Input_Signal,
       even2_Result(39) => Dangling_Input_Signal,
       even2_Result(40) => Dangling_Input_Signal,
       even2_Result(41) => Dangling_Input_Signal,
       even2_Result(42) => Dangling_Input_Signal,
       even2_Result(43) => Dangling_Input_Signal,
       even2_Result(44) => Dangling_Input_Signal,
       even2_Result(45) => Dangling_Input_Signal,
       even2_Result(46) => Dangling_Input_Signal,
       even2_Result(47) => Dangling_Input_Signal,
       even2_Result(48) => Dangling_Input_Signal,
       even2_Result(49) => Dangling_Input_Signal,
       even2_Result(50) => Dangling_Input_Signal,
       even2_Result(51) => Dangling_Input_Signal,
       even2_Result(52) => Dangling_Input_Signal,
       even2_Result(53) => Dangling_Input_Signal,
       even2_Result(54) => Dangling_Input_Signal,
       even2_Result(55) => Dangling_Input_Signal,
       even2_Result(56) => Dangling_Input_Signal,
       even2_Result(57) => Dangling_Input_Signal,
       even2_Result(58) => Dangling_Input_Signal,
       even2_Result(59) => Dangling_Input_Signal,
       even2_Result(60) => Dangling_Input_Signal,
       even2_Result(61) => Dangling_Input_Signal,
       even2_Result(62) => Dangling_Input_Signal,
       even2_Result(63) => Dangling_Input_Signal,
       even2_Result(64) => Dangling_Input_Signal,
       even2_Result(65) => Dangling_Input_Signal,
       even2_Result(66) => Dangling_Input_Signal,
       even2_Result(67) => Dangling_Input_Signal,
       even2_Result(68) => Dangling_Input_Signal,
       even2_Result(69) => Dangling_Input_Signal,
       even2_Result(70) => Dangling_Input_Signal,
       even2_Result(71) => Dangling_Input_Signal,
       even2_Result(72) => Dangling_Input_Signal,
       even2_Result(73) => Dangling_Input_Signal,
       even2_Result(74) => Dangling_Input_Signal,
       even2_Result(75) => Dangling_Input_Signal,
       even2_Result(76) => Dangling_Input_Signal,
       even2_Result(77) => Dangling_Input_Signal,
       even2_Result(78) => Dangling_Input_Signal,
       even2_Result(79) => Dangling_Input_Signal,
       even2_Result(80) => Dangling_Input_Signal,
       even2_Result(81) => Dangling_Input_Signal,
       even2_Result(82) => Dangling_Input_Signal,
       even2_Result(83) => Dangling_Input_Signal,
       even2_Result(84) => Dangling_Input_Signal,
       even2_Result(85) => Dangling_Input_Signal,
       even2_Result(86) => Dangling_Input_Signal,
       even2_Result(87) => Dangling_Input_Signal,
       even2_Result(88) => Dangling_Input_Signal,
       even2_Result(89) => Dangling_Input_Signal,
       even2_Result(90) => Dangling_Input_Signal,
       even2_Result(91) => Dangling_Input_Signal,
       even2_Result(92) => Dangling_Input_Signal,
       even2_Result(93) => Dangling_Input_Signal,
       even2_Result(94) => Dangling_Input_Signal,
       even2_Result(95) => Dangling_Input_Signal,
       even2_Result(96) => Dangling_Input_Signal,
       even2_Result(97) => Dangling_Input_Signal,
       even2_Result(98) => Dangling_Input_Signal,
       even2_Result(99) => Dangling_Input_Signal,
       even2_Result(100) => Dangling_Input_Signal,
       even2_Result(101) => Dangling_Input_Signal,
       even2_Result(102) => Dangling_Input_Signal,
       even2_Result(103) => Dangling_Input_Signal,
       even2_Result(104) => Dangling_Input_Signal,
       even2_Result(105) => Dangling_Input_Signal,
       even2_Result(106) => Dangling_Input_Signal,
       even2_Result(107) => Dangling_Input_Signal,
       even2_Result(108) => Dangling_Input_Signal,
       even2_Result(109) => Dangling_Input_Signal,
       even2_Result(110) => Dangling_Input_Signal,
       even2_Result(111) => Dangling_Input_Signal,
       even2_Result(112) => Dangling_Input_Signal,
       even2_Result(113) => Dangling_Input_Signal,
       even2_Result(114) => Dangling_Input_Signal,
       even2_Result(115) => Dangling_Input_Signal,
       even2_Result(116) => Dangling_Input_Signal,
       even2_Result(117) => Dangling_Input_Signal,
       even2_Result(118) => Dangling_Input_Signal,
       even2_Result(119) => Dangling_Input_Signal,
       even2_Result(120) => Dangling_Input_Signal,
       even2_Result(121) => Dangling_Input_Signal,
       even2_Result(122) => Dangling_Input_Signal,
       even2_Result(123) => Dangling_Input_Signal,
       even2_Result(124) => Dangling_Input_Signal,
       even2_Result(125) => Dangling_Input_Signal,
       even2_Result(126) => Dangling_Input_Signal,
       even2_Result(127) => Dangling_Input_Signal,
       even3_Latency(0) => Dangling_Input_Signal,
       even3_Latency(1) => Dangling_Input_Signal,
       even3_Latency(2) => Dangling_Input_Signal,
       even3_RegDst(0) => Dangling_Input_Signal,
       even3_RegDst(1) => Dangling_Input_Signal,
       even3_RegDst(2) => Dangling_Input_Signal,
       even3_RegDst(3) => Dangling_Input_Signal,
       even3_RegDst(4) => Dangling_Input_Signal,
       even3_RegDst(5) => Dangling_Input_Signal,
       even3_RegDst(6) => Dangling_Input_Signal,
       even3_Result(0) => Dangling_Input_Signal,
       even3_Result(1) => Dangling_Input_Signal,
       even3_Result(2) => Dangling_Input_Signal,
       even3_Result(3) => Dangling_Input_Signal,
       even3_Result(4) => Dangling_Input_Signal,
       even3_Result(5) => Dangling_Input_Signal,
       even3_Result(6) => Dangling_Input_Signal,
       even3_Result(7) => Dangling_Input_Signal,
       even3_Result(8) => Dangling_Input_Signal,
       even3_Result(9) => Dangling_Input_Signal,
       even3_Result(10) => Dangling_Input_Signal,
       even3_Result(11) => Dangling_Input_Signal,
       even3_Result(12) => Dangling_Input_Signal,
       even3_Result(13) => Dangling_Input_Signal,
       even3_Result(14) => Dangling_Input_Signal,
       even3_Result(15) => Dangling_Input_Signal,
       even3_Result(16) => Dangling_Input_Signal,
       even3_Result(17) => Dangling_Input_Signal,
       even3_Result(18) => Dangling_Input_Signal,
       even3_Result(19) => Dangling_Input_Signal,
       even3_Result(20) => Dangling_Input_Signal,
       even3_Result(21) => Dangling_Input_Signal,
       even3_Result(22) => Dangling_Input_Signal,
       even3_Result(23) => Dangling_Input_Signal,
       even3_Result(24) => Dangling_Input_Signal,
       even3_Result(25) => Dangling_Input_Signal,
       even3_Result(26) => Dangling_Input_Signal,
       even3_Result(27) => Dangling_Input_Signal,
       even3_Result(28) => Dangling_Input_Signal,
       even3_Result(29) => Dangling_Input_Signal,
       even3_Result(30) => Dangling_Input_Signal,
       even3_Result(31) => Dangling_Input_Signal,
       even3_Result(32) => Dangling_Input_Signal,
       even3_Result(33) => Dangling_Input_Signal,
       even3_Result(34) => Dangling_Input_Signal,
       even3_Result(35) => Dangling_Input_Signal,
       even3_Result(36) => Dangling_Input_Signal,
       even3_Result(37) => Dangling_Input_Signal,
       even3_Result(38) => Dangling_Input_Signal,
       even3_Result(39) => Dangling_Input_Signal,
       even3_Result(40) => Dangling_Input_Signal,
       even3_Result(41) => Dangling_Input_Signal,
       even3_Result(42) => Dangling_Input_Signal,
       even3_Result(43) => Dangling_Input_Signal,
       even3_Result(44) => Dangling_Input_Signal,
       even3_Result(45) => Dangling_Input_Signal,
       even3_Result(46) => Dangling_Input_Signal,
       even3_Result(47) => Dangling_Input_Signal,
       even3_Result(48) => Dangling_Input_Signal,
       even3_Result(49) => Dangling_Input_Signal,
       even3_Result(50) => Dangling_Input_Signal,
       even3_Result(51) => Dangling_Input_Signal,
       even3_Result(52) => Dangling_Input_Signal,
       even3_Result(53) => Dangling_Input_Signal,
       even3_Result(54) => Dangling_Input_Signal,
       even3_Result(55) => Dangling_Input_Signal,
       even3_Result(56) => Dangling_Input_Signal,
       even3_Result(57) => Dangling_Input_Signal,
       even3_Result(58) => Dangling_Input_Signal,
       even3_Result(59) => Dangling_Input_Signal,
       even3_Result(60) => Dangling_Input_Signal,
       even3_Result(61) => Dangling_Input_Signal,
       even3_Result(62) => Dangling_Input_Signal,
       even3_Result(63) => Dangling_Input_Signal,
       even3_Result(64) => Dangling_Input_Signal,
       even3_Result(65) => Dangling_Input_Signal,
       even3_Result(66) => Dangling_Input_Signal,
       even3_Result(67) => Dangling_Input_Signal,
       even3_Result(68) => Dangling_Input_Signal,
       even3_Result(69) => Dangling_Input_Signal,
       even3_Result(70) => Dangling_Input_Signal,
       even3_Result(71) => Dangling_Input_Signal,
       even3_Result(72) => Dangling_Input_Signal,
       even3_Result(73) => Dangling_Input_Signal,
       even3_Result(74) => Dangling_Input_Signal,
       even3_Result(75) => Dangling_Input_Signal,
       even3_Result(76) => Dangling_Input_Signal,
       even3_Result(77) => Dangling_Input_Signal,
       even3_Result(78) => Dangling_Input_Signal,
       even3_Result(79) => Dangling_Input_Signal,
       even3_Result(80) => Dangling_Input_Signal,
       even3_Result(81) => Dangling_Input_Signal,
       even3_Result(82) => Dangling_Input_Signal,
       even3_Result(83) => Dangling_Input_Signal,
       even3_Result(84) => Dangling_Input_Signal,
       even3_Result(85) => Dangling_Input_Signal,
       even3_Result(86) => Dangling_Input_Signal,
       even3_Result(87) => Dangling_Input_Signal,
       even3_Result(88) => Dangling_Input_Signal,
       even3_Result(89) => Dangling_Input_Signal,
       even3_Result(90) => Dangling_Input_Signal,
       even3_Result(91) => Dangling_Input_Signal,
       even3_Result(92) => Dangling_Input_Signal,
       even3_Result(93) => Dangling_Input_Signal,
       even3_Result(94) => Dangling_Input_Signal,
       even3_Result(95) => Dangling_Input_Signal,
       even3_Result(96) => Dangling_Input_Signal,
       even3_Result(97) => Dangling_Input_Signal,
       even3_Result(98) => Dangling_Input_Signal,
       even3_Result(99) => Dangling_Input_Signal,
       even3_Result(100) => Dangling_Input_Signal,
       even3_Result(101) => Dangling_Input_Signal,
       even3_Result(102) => Dangling_Input_Signal,
       even3_Result(103) => Dangling_Input_Signal,
       even3_Result(104) => Dangling_Input_Signal,
       even3_Result(105) => Dangling_Input_Signal,
       even3_Result(106) => Dangling_Input_Signal,
       even3_Result(107) => Dangling_Input_Signal,
       even3_Result(108) => Dangling_Input_Signal,
       even3_Result(109) => Dangling_Input_Signal,
       even3_Result(110) => Dangling_Input_Signal,
       even3_Result(111) => Dangling_Input_Signal,
       even3_Result(112) => Dangling_Input_Signal,
       even3_Result(113) => Dangling_Input_Signal,
       even3_Result(114) => Dangling_Input_Signal,
       even3_Result(115) => Dangling_Input_Signal,
       even3_Result(116) => Dangling_Input_Signal,
       even3_Result(117) => Dangling_Input_Signal,
       even3_Result(118) => Dangling_Input_Signal,
       even3_Result(119) => Dangling_Input_Signal,
       even3_Result(120) => Dangling_Input_Signal,
       even3_Result(121) => Dangling_Input_Signal,
       even3_Result(122) => Dangling_Input_Signal,
       even3_Result(123) => Dangling_Input_Signal,
       even3_Result(124) => Dangling_Input_Signal,
       even3_Result(125) => Dangling_Input_Signal,
       even3_Result(126) => Dangling_Input_Signal,
       even3_Result(127) => Dangling_Input_Signal,
       even4_Latency(0) => Dangling_Input_Signal,
       even4_Latency(1) => Dangling_Input_Signal,
       even4_Latency(2) => Dangling_Input_Signal,
       even4_RegDst(0) => Dangling_Input_Signal,
       even4_RegDst(1) => Dangling_Input_Signal,
       even4_RegDst(2) => Dangling_Input_Signal,
       even4_RegDst(3) => Dangling_Input_Signal,
       even4_RegDst(4) => Dangling_Input_Signal,
       even4_RegDst(5) => Dangling_Input_Signal,
       even4_RegDst(6) => Dangling_Input_Signal,
       even4_Result(0) => Dangling_Input_Signal,
       even4_Result(1) => Dangling_Input_Signal,
       even4_Result(2) => Dangling_Input_Signal,
       even4_Result(3) => Dangling_Input_Signal,
       even4_Result(4) => Dangling_Input_Signal,
       even4_Result(5) => Dangling_Input_Signal,
       even4_Result(6) => Dangling_Input_Signal,
       even4_Result(7) => Dangling_Input_Signal,
       even4_Result(8) => Dangling_Input_Signal,
       even4_Result(9) => Dangling_Input_Signal,
       even4_Result(10) => Dangling_Input_Signal,
       even4_Result(11) => Dangling_Input_Signal,
       even4_Result(12) => Dangling_Input_Signal,
       even4_Result(13) => Dangling_Input_Signal,
       even4_Result(14) => Dangling_Input_Signal,
       even4_Result(15) => Dangling_Input_Signal,
       even4_Result(16) => Dangling_Input_Signal,
       even4_Result(17) => Dangling_Input_Signal,
       even4_Result(18) => Dangling_Input_Signal,
       even4_Result(19) => Dangling_Input_Signal,
       even4_Result(20) => Dangling_Input_Signal,
       even4_Result(21) => Dangling_Input_Signal,
       even4_Result(22) => Dangling_Input_Signal,
       even4_Result(23) => Dangling_Input_Signal,
       even4_Result(24) => Dangling_Input_Signal,
       even4_Result(25) => Dangling_Input_Signal,
       even4_Result(26) => Dangling_Input_Signal,
       even4_Result(27) => Dangling_Input_Signal,
       even4_Result(28) => Dangling_Input_Signal,
       even4_Result(29) => Dangling_Input_Signal,
       even4_Result(30) => Dangling_Input_Signal,
       even4_Result(31) => Dangling_Input_Signal,
       even4_Result(32) => Dangling_Input_Signal,
       even4_Result(33) => Dangling_Input_Signal,
       even4_Result(34) => Dangling_Input_Signal,
       even4_Result(35) => Dangling_Input_Signal,
       even4_Result(36) => Dangling_Input_Signal,
       even4_Result(37) => Dangling_Input_Signal,
       even4_Result(38) => Dangling_Input_Signal,
       even4_Result(39) => Dangling_Input_Signal,
       even4_Result(40) => Dangling_Input_Signal,
       even4_Result(41) => Dangling_Input_Signal,
       even4_Result(42) => Dangling_Input_Signal,
       even4_Result(43) => Dangling_Input_Signal,
       even4_Result(44) => Dangling_Input_Signal,
       even4_Result(45) => Dangling_Input_Signal,
       even4_Result(46) => Dangling_Input_Signal,
       even4_Result(47) => Dangling_Input_Signal,
       even4_Result(48) => Dangling_Input_Signal,
       even4_Result(49) => Dangling_Input_Signal,
       even4_Result(50) => Dangling_Input_Signal,
       even4_Result(51) => Dangling_Input_Signal,
       even4_Result(52) => Dangling_Input_Signal,
       even4_Result(53) => Dangling_Input_Signal,
       even4_Result(54) => Dangling_Input_Signal,
       even4_Result(55) => Dangling_Input_Signal,
       even4_Result(56) => Dangling_Input_Signal,
       even4_Result(57) => Dangling_Input_Signal,
       even4_Result(58) => Dangling_Input_Signal,
       even4_Result(59) => Dangling_Input_Signal,
       even4_Result(60) => Dangling_Input_Signal,
       even4_Result(61) => Dangling_Input_Signal,
       even4_Result(62) => Dangling_Input_Signal,
       even4_Result(63) => Dangling_Input_Signal,
       even4_Result(64) => Dangling_Input_Signal,
       even4_Result(65) => Dangling_Input_Signal,
       even4_Result(66) => Dangling_Input_Signal,
       even4_Result(67) => Dangling_Input_Signal,
       even4_Result(68) => Dangling_Input_Signal,
       even4_Result(69) => Dangling_Input_Signal,
       even4_Result(70) => Dangling_Input_Signal,
       even4_Result(71) => Dangling_Input_Signal,
       even4_Result(72) => Dangling_Input_Signal,
       even4_Result(73) => Dangling_Input_Signal,
       even4_Result(74) => Dangling_Input_Signal,
       even4_Result(75) => Dangling_Input_Signal,
       even4_Result(76) => Dangling_Input_Signal,
       even4_Result(77) => Dangling_Input_Signal,
       even4_Result(78) => Dangling_Input_Signal,
       even4_Result(79) => Dangling_Input_Signal,
       even4_Result(80) => Dangling_Input_Signal,
       even4_Result(81) => Dangling_Input_Signal,
       even4_Result(82) => Dangling_Input_Signal,
       even4_Result(83) => Dangling_Input_Signal,
       even4_Result(84) => Dangling_Input_Signal,
       even4_Result(85) => Dangling_Input_Signal,
       even4_Result(86) => Dangling_Input_Signal,
       even4_Result(87) => Dangling_Input_Signal,
       even4_Result(88) => Dangling_Input_Signal,
       even4_Result(89) => Dangling_Input_Signal,
       even4_Result(90) => Dangling_Input_Signal,
       even4_Result(91) => Dangling_Input_Signal,
       even4_Result(92) => Dangling_Input_Signal,
       even4_Result(93) => Dangling_Input_Signal,
       even4_Result(94) => Dangling_Input_Signal,
       even4_Result(95) => Dangling_Input_Signal,
       even4_Result(96) => Dangling_Input_Signal,
       even4_Result(97) => Dangling_Input_Signal,
       even4_Result(98) => Dangling_Input_Signal,
       even4_Result(99) => Dangling_Input_Signal,
       even4_Result(100) => Dangling_Input_Signal,
       even4_Result(101) => Dangling_Input_Signal,
       even4_Result(102) => Dangling_Input_Signal,
       even4_Result(103) => Dangling_Input_Signal,
       even4_Result(104) => Dangling_Input_Signal,
       even4_Result(105) => Dangling_Input_Signal,
       even4_Result(106) => Dangling_Input_Signal,
       even4_Result(107) => Dangling_Input_Signal,
       even4_Result(108) => Dangling_Input_Signal,
       even4_Result(109) => Dangling_Input_Signal,
       even4_Result(110) => Dangling_Input_Signal,
       even4_Result(111) => Dangling_Input_Signal,
       even4_Result(112) => Dangling_Input_Signal,
       even4_Result(113) => Dangling_Input_Signal,
       even4_Result(114) => Dangling_Input_Signal,
       even4_Result(115) => Dangling_Input_Signal,
       even4_Result(116) => Dangling_Input_Signal,
       even4_Result(117) => Dangling_Input_Signal,
       even4_Result(118) => Dangling_Input_Signal,
       even4_Result(119) => Dangling_Input_Signal,
       even4_Result(120) => Dangling_Input_Signal,
       even4_Result(121) => Dangling_Input_Signal,
       even4_Result(122) => Dangling_Input_Signal,
       even4_Result(123) => Dangling_Input_Signal,
       even4_Result(124) => Dangling_Input_Signal,
       even4_Result(125) => Dangling_Input_Signal,
       even4_Result(126) => Dangling_Input_Signal,
       even4_Result(127) => Dangling_Input_Signal,
       even5_Latency(0) => Dangling_Input_Signal,
       even5_Latency(1) => Dangling_Input_Signal,
       even5_Latency(2) => Dangling_Input_Signal,
       even5_RegDst(0) => Dangling_Input_Signal,
       even5_RegDst(1) => Dangling_Input_Signal,
       even5_RegDst(2) => Dangling_Input_Signal,
       even5_RegDst(3) => Dangling_Input_Signal,
       even5_RegDst(4) => Dangling_Input_Signal,
       even5_RegDst(5) => Dangling_Input_Signal,
       even5_RegDst(6) => Dangling_Input_Signal,
       even5_Result(0) => Dangling_Input_Signal,
       even5_Result(1) => Dangling_Input_Signal,
       even5_Result(2) => Dangling_Input_Signal,
       even5_Result(3) => Dangling_Input_Signal,
       even5_Result(4) => Dangling_Input_Signal,
       even5_Result(5) => Dangling_Input_Signal,
       even5_Result(6) => Dangling_Input_Signal,
       even5_Result(7) => Dangling_Input_Signal,
       even5_Result(8) => Dangling_Input_Signal,
       even5_Result(9) => Dangling_Input_Signal,
       even5_Result(10) => Dangling_Input_Signal,
       even5_Result(11) => Dangling_Input_Signal,
       even5_Result(12) => Dangling_Input_Signal,
       even5_Result(13) => Dangling_Input_Signal,
       even5_Result(14) => Dangling_Input_Signal,
       even5_Result(15) => Dangling_Input_Signal,
       even5_Result(16) => Dangling_Input_Signal,
       even5_Result(17) => Dangling_Input_Signal,
       even5_Result(18) => Dangling_Input_Signal,
       even5_Result(19) => Dangling_Input_Signal,
       even5_Result(20) => Dangling_Input_Signal,
       even5_Result(21) => Dangling_Input_Signal,
       even5_Result(22) => Dangling_Input_Signal,
       even5_Result(23) => Dangling_Input_Signal,
       even5_Result(24) => Dangling_Input_Signal,
       even5_Result(25) => Dangling_Input_Signal,
       even5_Result(26) => Dangling_Input_Signal,
       even5_Result(27) => Dangling_Input_Signal,
       even5_Result(28) => Dangling_Input_Signal,
       even5_Result(29) => Dangling_Input_Signal,
       even5_Result(30) => Dangling_Input_Signal,
       even5_Result(31) => Dangling_Input_Signal,
       even5_Result(32) => Dangling_Input_Signal,
       even5_Result(33) => Dangling_Input_Signal,
       even5_Result(34) => Dangling_Input_Signal,
       even5_Result(35) => Dangling_Input_Signal,
       even5_Result(36) => Dangling_Input_Signal,
       even5_Result(37) => Dangling_Input_Signal,
       even5_Result(38) => Dangling_Input_Signal,
       even5_Result(39) => Dangling_Input_Signal,
       even5_Result(40) => Dangling_Input_Signal,
       even5_Result(41) => Dangling_Input_Signal,
       even5_Result(42) => Dangling_Input_Signal,
       even5_Result(43) => Dangling_Input_Signal,
       even5_Result(44) => Dangling_Input_Signal,
       even5_Result(45) => Dangling_Input_Signal,
       even5_Result(46) => Dangling_Input_Signal,
       even5_Result(47) => Dangling_Input_Signal,
       even5_Result(48) => Dangling_Input_Signal,
       even5_Result(49) => Dangling_Input_Signal,
       even5_Result(50) => Dangling_Input_Signal,
       even5_Result(51) => Dangling_Input_Signal,
       even5_Result(52) => Dangling_Input_Signal,
       even5_Result(53) => Dangling_Input_Signal,
       even5_Result(54) => Dangling_Input_Signal,
       even5_Result(55) => Dangling_Input_Signal,
       even5_Result(56) => Dangling_Input_Signal,
       even5_Result(57) => Dangling_Input_Signal,
       even5_Result(58) => Dangling_Input_Signal,
       even5_Result(59) => Dangling_Input_Signal,
       even5_Result(60) => Dangling_Input_Signal,
       even5_Result(61) => Dangling_Input_Signal,
       even5_Result(62) => Dangling_Input_Signal,
       even5_Result(63) => Dangling_Input_Signal,
       even5_Result(64) => Dangling_Input_Signal,
       even5_Result(65) => Dangling_Input_Signal,
       even5_Result(66) => Dangling_Input_Signal,
       even5_Result(67) => Dangling_Input_Signal,
       even5_Result(68) => Dangling_Input_Signal,
       even5_Result(69) => Dangling_Input_Signal,
       even5_Result(70) => Dangling_Input_Signal,
       even5_Result(71) => Dangling_Input_Signal,
       even5_Result(72) => Dangling_Input_Signal,
       even5_Result(73) => Dangling_Input_Signal,
       even5_Result(74) => Dangling_Input_Signal,
       even5_Result(75) => Dangling_Input_Signal,
       even5_Result(76) => Dangling_Input_Signal,
       even5_Result(77) => Dangling_Input_Signal,
       even5_Result(78) => Dangling_Input_Signal,
       even5_Result(79) => Dangling_Input_Signal,
       even5_Result(80) => Dangling_Input_Signal,
       even5_Result(81) => Dangling_Input_Signal,
       even5_Result(82) => Dangling_Input_Signal,
       even5_Result(83) => Dangling_Input_Signal,
       even5_Result(84) => Dangling_Input_Signal,
       even5_Result(85) => Dangling_Input_Signal,
       even5_Result(86) => Dangling_Input_Signal,
       even5_Result(87) => Dangling_Input_Signal,
       even5_Result(88) => Dangling_Input_Signal,
       even5_Result(89) => Dangling_Input_Signal,
       even5_Result(90) => Dangling_Input_Signal,
       even5_Result(91) => Dangling_Input_Signal,
       even5_Result(92) => Dangling_Input_Signal,
       even5_Result(93) => Dangling_Input_Signal,
       even5_Result(94) => Dangling_Input_Signal,
       even5_Result(95) => Dangling_Input_Signal,
       even5_Result(96) => Dangling_Input_Signal,
       even5_Result(97) => Dangling_Input_Signal,
       even5_Result(98) => Dangling_Input_Signal,
       even5_Result(99) => Dangling_Input_Signal,
       even5_Result(100) => Dangling_Input_Signal,
       even5_Result(101) => Dangling_Input_Signal,
       even5_Result(102) => Dangling_Input_Signal,
       even5_Result(103) => Dangling_Input_Signal,
       even5_Result(104) => Dangling_Input_Signal,
       even5_Result(105) => Dangling_Input_Signal,
       even5_Result(106) => Dangling_Input_Signal,
       even5_Result(107) => Dangling_Input_Signal,
       even5_Result(108) => Dangling_Input_Signal,
       even5_Result(109) => Dangling_Input_Signal,
       even5_Result(110) => Dangling_Input_Signal,
       even5_Result(111) => Dangling_Input_Signal,
       even5_Result(112) => Dangling_Input_Signal,
       even5_Result(113) => Dangling_Input_Signal,
       even5_Result(114) => Dangling_Input_Signal,
       even5_Result(115) => Dangling_Input_Signal,
       even5_Result(116) => Dangling_Input_Signal,
       even5_Result(117) => Dangling_Input_Signal,
       even5_Result(118) => Dangling_Input_Signal,
       even5_Result(119) => Dangling_Input_Signal,
       even5_Result(120) => Dangling_Input_Signal,
       even5_Result(121) => Dangling_Input_Signal,
       even5_Result(122) => Dangling_Input_Signal,
       even5_Result(123) => Dangling_Input_Signal,
       even5_Result(124) => Dangling_Input_Signal,
       even5_Result(125) => Dangling_Input_Signal,
       even5_Result(126) => Dangling_Input_Signal,
       even5_Result(127) => Dangling_Input_Signal,
       even6_Latency(0) => Dangling_Input_Signal,
       even6_Latency(1) => Dangling_Input_Signal,
       even6_Latency(2) => Dangling_Input_Signal,
       even6_RegDst(0) => Dangling_Input_Signal,
       even6_RegDst(1) => Dangling_Input_Signal,
       even6_RegDst(2) => Dangling_Input_Signal,
       even6_RegDst(3) => Dangling_Input_Signal,
       even6_RegDst(4) => Dangling_Input_Signal,
       even6_RegDst(5) => Dangling_Input_Signal,
       even6_RegDst(6) => Dangling_Input_Signal,
       even6_Result(0) => Dangling_Input_Signal,
       even6_Result(1) => Dangling_Input_Signal,
       even6_Result(2) => Dangling_Input_Signal,
       even6_Result(3) => Dangling_Input_Signal,
       even6_Result(4) => Dangling_Input_Signal,
       even6_Result(5) => Dangling_Input_Signal,
       even6_Result(6) => Dangling_Input_Signal,
       even6_Result(7) => Dangling_Input_Signal,
       even6_Result(8) => Dangling_Input_Signal,
       even6_Result(9) => Dangling_Input_Signal,
       even6_Result(10) => Dangling_Input_Signal,
       even6_Result(11) => Dangling_Input_Signal,
       even6_Result(12) => Dangling_Input_Signal,
       even6_Result(13) => Dangling_Input_Signal,
       even6_Result(14) => Dangling_Input_Signal,
       even6_Result(15) => Dangling_Input_Signal,
       even6_Result(16) => Dangling_Input_Signal,
       even6_Result(17) => Dangling_Input_Signal,
       even6_Result(18) => Dangling_Input_Signal,
       even6_Result(19) => Dangling_Input_Signal,
       even6_Result(20) => Dangling_Input_Signal,
       even6_Result(21) => Dangling_Input_Signal,
       even6_Result(22) => Dangling_Input_Signal,
       even6_Result(23) => Dangling_Input_Signal,
       even6_Result(24) => Dangling_Input_Signal,
       even6_Result(25) => Dangling_Input_Signal,
       even6_Result(26) => Dangling_Input_Signal,
       even6_Result(27) => Dangling_Input_Signal,
       even6_Result(28) => Dangling_Input_Signal,
       even6_Result(29) => Dangling_Input_Signal,
       even6_Result(30) => Dangling_Input_Signal,
       even6_Result(31) => Dangling_Input_Signal,
       even6_Result(32) => Dangling_Input_Signal,
       even6_Result(33) => Dangling_Input_Signal,
       even6_Result(34) => Dangling_Input_Signal,
       even6_Result(35) => Dangling_Input_Signal,
       even6_Result(36) => Dangling_Input_Signal,
       even6_Result(37) => Dangling_Input_Signal,
       even6_Result(38) => Dangling_Input_Signal,
       even6_Result(39) => Dangling_Input_Signal,
       even6_Result(40) => Dangling_Input_Signal,
       even6_Result(41) => Dangling_Input_Signal,
       even6_Result(42) => Dangling_Input_Signal,
       even6_Result(43) => Dangling_Input_Signal,
       even6_Result(44) => Dangling_Input_Signal,
       even6_Result(45) => Dangling_Input_Signal,
       even6_Result(46) => Dangling_Input_Signal,
       even6_Result(47) => Dangling_Input_Signal,
       even6_Result(48) => Dangling_Input_Signal,
       even6_Result(49) => Dangling_Input_Signal,
       even6_Result(50) => Dangling_Input_Signal,
       even6_Result(51) => Dangling_Input_Signal,
       even6_Result(52) => Dangling_Input_Signal,
       even6_Result(53) => Dangling_Input_Signal,
       even6_Result(54) => Dangling_Input_Signal,
       even6_Result(55) => Dangling_Input_Signal,
       even6_Result(56) => Dangling_Input_Signal,
       even6_Result(57) => Dangling_Input_Signal,
       even6_Result(58) => Dangling_Input_Signal,
       even6_Result(59) => Dangling_Input_Signal,
       even6_Result(60) => Dangling_Input_Signal,
       even6_Result(61) => Dangling_Input_Signal,
       even6_Result(62) => Dangling_Input_Signal,
       even6_Result(63) => Dangling_Input_Signal,
       even6_Result(64) => Dangling_Input_Signal,
       even6_Result(65) => Dangling_Input_Signal,
       even6_Result(66) => Dangling_Input_Signal,
       even6_Result(67) => Dangling_Input_Signal,
       even6_Result(68) => Dangling_Input_Signal,
       even6_Result(69) => Dangling_Input_Signal,
       even6_Result(70) => Dangling_Input_Signal,
       even6_Result(71) => Dangling_Input_Signal,
       even6_Result(72) => Dangling_Input_Signal,
       even6_Result(73) => Dangling_Input_Signal,
       even6_Result(74) => Dangling_Input_Signal,
       even6_Result(75) => Dangling_Input_Signal,
       even6_Result(76) => Dangling_Input_Signal,
       even6_Result(77) => Dangling_Input_Signal,
       even6_Result(78) => Dangling_Input_Signal,
       even6_Result(79) => Dangling_Input_Signal,
       even6_Result(80) => Dangling_Input_Signal,
       even6_Result(81) => Dangling_Input_Signal,
       even6_Result(82) => Dangling_Input_Signal,
       even6_Result(83) => Dangling_Input_Signal,
       even6_Result(84) => Dangling_Input_Signal,
       even6_Result(85) => Dangling_Input_Signal,
       even6_Result(86) => Dangling_Input_Signal,
       even6_Result(87) => Dangling_Input_Signal,
       even6_Result(88) => Dangling_Input_Signal,
       even6_Result(89) => Dangling_Input_Signal,
       even6_Result(90) => Dangling_Input_Signal,
       even6_Result(91) => Dangling_Input_Signal,
       even6_Result(92) => Dangling_Input_Signal,
       even6_Result(93) => Dangling_Input_Signal,
       even6_Result(94) => Dangling_Input_Signal,
       even6_Result(95) => Dangling_Input_Signal,
       even6_Result(96) => Dangling_Input_Signal,
       even6_Result(97) => Dangling_Input_Signal,
       even6_Result(98) => Dangling_Input_Signal,
       even6_Result(99) => Dangling_Input_Signal,
       even6_Result(100) => Dangling_Input_Signal,
       even6_Result(101) => Dangling_Input_Signal,
       even6_Result(102) => Dangling_Input_Signal,
       even6_Result(103) => Dangling_Input_Signal,
       even6_Result(104) => Dangling_Input_Signal,
       even6_Result(105) => Dangling_Input_Signal,
       even6_Result(106) => Dangling_Input_Signal,
       even6_Result(107) => Dangling_Input_Signal,
       even6_Result(108) => Dangling_Input_Signal,
       even6_Result(109) => Dangling_Input_Signal,
       even6_Result(110) => Dangling_Input_Signal,
       even6_Result(111) => Dangling_Input_Signal,
       even6_Result(112) => Dangling_Input_Signal,
       even6_Result(113) => Dangling_Input_Signal,
       even6_Result(114) => Dangling_Input_Signal,
       even6_Result(115) => Dangling_Input_Signal,
       even6_Result(116) => Dangling_Input_Signal,
       even6_Result(117) => Dangling_Input_Signal,
       even6_Result(118) => Dangling_Input_Signal,
       even6_Result(119) => Dangling_Input_Signal,
       even6_Result(120) => Dangling_Input_Signal,
       even6_Result(121) => Dangling_Input_Signal,
       even6_Result(122) => Dangling_Input_Signal,
       even6_Result(123) => Dangling_Input_Signal,
       even6_Result(124) => Dangling_Input_Signal,
       even6_Result(125) => Dangling_Input_Signal,
       even6_Result(126) => Dangling_Input_Signal,
       even6_Result(127) => Dangling_Input_Signal,
       even7_Latency(0) => Dangling_Input_Signal,
       even7_Latency(1) => Dangling_Input_Signal,
       even7_Latency(2) => Dangling_Input_Signal,
       even7_RegDst(0) => Dangling_Input_Signal,
       even7_RegDst(1) => Dangling_Input_Signal,
       even7_RegDst(2) => Dangling_Input_Signal,
       even7_RegDst(3) => Dangling_Input_Signal,
       even7_RegDst(4) => Dangling_Input_Signal,
       even7_RegDst(5) => Dangling_Input_Signal,
       even7_RegDst(6) => Dangling_Input_Signal,
       even7_Result(0) => Dangling_Input_Signal,
       even7_Result(1) => Dangling_Input_Signal,
       even7_Result(2) => Dangling_Input_Signal,
       even7_Result(3) => Dangling_Input_Signal,
       even7_Result(4) => Dangling_Input_Signal,
       even7_Result(5) => Dangling_Input_Signal,
       even7_Result(6) => Dangling_Input_Signal,
       even7_Result(7) => Dangling_Input_Signal,
       even7_Result(8) => Dangling_Input_Signal,
       even7_Result(9) => Dangling_Input_Signal,
       even7_Result(10) => Dangling_Input_Signal,
       even7_Result(11) => Dangling_Input_Signal,
       even7_Result(12) => Dangling_Input_Signal,
       even7_Result(13) => Dangling_Input_Signal,
       even7_Result(14) => Dangling_Input_Signal,
       even7_Result(15) => Dangling_Input_Signal,
       even7_Result(16) => Dangling_Input_Signal,
       even7_Result(17) => Dangling_Input_Signal,
       even7_Result(18) => Dangling_Input_Signal,
       even7_Result(19) => Dangling_Input_Signal,
       even7_Result(20) => Dangling_Input_Signal,
       even7_Result(21) => Dangling_Input_Signal,
       even7_Result(22) => Dangling_Input_Signal,
       even7_Result(23) => Dangling_Input_Signal,
       even7_Result(24) => Dangling_Input_Signal,
       even7_Result(25) => Dangling_Input_Signal,
       even7_Result(26) => Dangling_Input_Signal,
       even7_Result(27) => Dangling_Input_Signal,
       even7_Result(28) => Dangling_Input_Signal,
       even7_Result(29) => Dangling_Input_Signal,
       even7_Result(30) => Dangling_Input_Signal,
       even7_Result(31) => Dangling_Input_Signal,
       even7_Result(32) => Dangling_Input_Signal,
       even7_Result(33) => Dangling_Input_Signal,
       even7_Result(34) => Dangling_Input_Signal,
       even7_Result(35) => Dangling_Input_Signal,
       even7_Result(36) => Dangling_Input_Signal,
       even7_Result(37) => Dangling_Input_Signal,
       even7_Result(38) => Dangling_Input_Signal,
       even7_Result(39) => Dangling_Input_Signal,
       even7_Result(40) => Dangling_Input_Signal,
       even7_Result(41) => Dangling_Input_Signal,
       even7_Result(42) => Dangling_Input_Signal,
       even7_Result(43) => Dangling_Input_Signal,
       even7_Result(44) => Dangling_Input_Signal,
       even7_Result(45) => Dangling_Input_Signal,
       even7_Result(46) => Dangling_Input_Signal,
       even7_Result(47) => Dangling_Input_Signal,
       even7_Result(48) => Dangling_Input_Signal,
       even7_Result(49) => Dangling_Input_Signal,
       even7_Result(50) => Dangling_Input_Signal,
       even7_Result(51) => Dangling_Input_Signal,
       even7_Result(52) => Dangling_Input_Signal,
       even7_Result(53) => Dangling_Input_Signal,
       even7_Result(54) => Dangling_Input_Signal,
       even7_Result(55) => Dangling_Input_Signal,
       even7_Result(56) => Dangling_Input_Signal,
       even7_Result(57) => Dangling_Input_Signal,
       even7_Result(58) => Dangling_Input_Signal,
       even7_Result(59) => Dangling_Input_Signal,
       even7_Result(60) => Dangling_Input_Signal,
       even7_Result(61) => Dangling_Input_Signal,
       even7_Result(62) => Dangling_Input_Signal,
       even7_Result(63) => Dangling_Input_Signal,
       even7_Result(64) => Dangling_Input_Signal,
       even7_Result(65) => Dangling_Input_Signal,
       even7_Result(66) => Dangling_Input_Signal,
       even7_Result(67) => Dangling_Input_Signal,
       even7_Result(68) => Dangling_Input_Signal,
       even7_Result(69) => Dangling_Input_Signal,
       even7_Result(70) => Dangling_Input_Signal,
       even7_Result(71) => Dangling_Input_Signal,
       even7_Result(72) => Dangling_Input_Signal,
       even7_Result(73) => Dangling_Input_Signal,
       even7_Result(74) => Dangling_Input_Signal,
       even7_Result(75) => Dangling_Input_Signal,
       even7_Result(76) => Dangling_Input_Signal,
       even7_Result(77) => Dangling_Input_Signal,
       even7_Result(78) => Dangling_Input_Signal,
       even7_Result(79) => Dangling_Input_Signal,
       even7_Result(80) => Dangling_Input_Signal,
       even7_Result(81) => Dangling_Input_Signal,
       even7_Result(82) => Dangling_Input_Signal,
       even7_Result(83) => Dangling_Input_Signal,
       even7_Result(84) => Dangling_Input_Signal,
       even7_Result(85) => Dangling_Input_Signal,
       even7_Result(86) => Dangling_Input_Signal,
       even7_Result(87) => Dangling_Input_Signal,
       even7_Result(88) => Dangling_Input_Signal,
       even7_Result(89) => Dangling_Input_Signal,
       even7_Result(90) => Dangling_Input_Signal,
       even7_Result(91) => Dangling_Input_Signal,
       even7_Result(92) => Dangling_Input_Signal,
       even7_Result(93) => Dangling_Input_Signal,
       even7_Result(94) => Dangling_Input_Signal,
       even7_Result(95) => Dangling_Input_Signal,
       even7_Result(96) => Dangling_Input_Signal,
       even7_Result(97) => Dangling_Input_Signal,
       even7_Result(98) => Dangling_Input_Signal,
       even7_Result(99) => Dangling_Input_Signal,
       even7_Result(100) => Dangling_Input_Signal,
       even7_Result(101) => Dangling_Input_Signal,
       even7_Result(102) => Dangling_Input_Signal,
       even7_Result(103) => Dangling_Input_Signal,
       even7_Result(104) => Dangling_Input_Signal,
       even7_Result(105) => Dangling_Input_Signal,
       even7_Result(106) => Dangling_Input_Signal,
       even7_Result(107) => Dangling_Input_Signal,
       even7_Result(108) => Dangling_Input_Signal,
       even7_Result(109) => Dangling_Input_Signal,
       even7_Result(110) => Dangling_Input_Signal,
       even7_Result(111) => Dangling_Input_Signal,
       even7_Result(112) => Dangling_Input_Signal,
       even7_Result(113) => Dangling_Input_Signal,
       even7_Result(114) => Dangling_Input_Signal,
       even7_Result(115) => Dangling_Input_Signal,
       even7_Result(116) => Dangling_Input_Signal,
       even7_Result(117) => Dangling_Input_Signal,
       even7_Result(118) => Dangling_Input_Signal,
       even7_Result(119) => Dangling_Input_Signal,
       even7_Result(120) => Dangling_Input_Signal,
       even7_Result(121) => Dangling_Input_Signal,
       even7_Result(122) => Dangling_Input_Signal,
       even7_Result(123) => Dangling_Input_Signal,
       even7_Result(124) => Dangling_Input_Signal,
       even7_Result(125) => Dangling_Input_Signal,
       even7_Result(126) => Dangling_Input_Signal,
       even7_Result(127) => Dangling_Input_Signal,
       E_reg(0) => Dangling_Input_Signal,
       E_reg(1) => Dangling_Input_Signal,
       E_reg(2) => Dangling_Input_Signal,
       E_reg(3) => Dangling_Input_Signal,
       E_reg(4) => Dangling_Input_Signal,
       E_reg(5) => Dangling_Input_Signal,
       E_reg(6) => Dangling_Input_Signal,
       E_reg(7) => Dangling_Input_Signal,
       E_reg(8) => Dangling_Input_Signal,
       E_reg(9) => Dangling_Input_Signal,
       E_reg(10) => Dangling_Input_Signal,
       E_reg(11) => Dangling_Input_Signal,
       E_reg(12) => Dangling_Input_Signal,
       E_reg(13) => Dangling_Input_Signal,
       E_reg(14) => Dangling_Input_Signal,
       E_reg(15) => Dangling_Input_Signal,
       E_reg(16) => Dangling_Input_Signal,
       E_reg(17) => Dangling_Input_Signal,
       E_reg(18) => Dangling_Input_Signal,
       E_reg(19) => Dangling_Input_Signal,
       E_reg(20) => Dangling_Input_Signal,
       E_reg(21) => Dangling_Input_Signal,
       E_reg(22) => Dangling_Input_Signal,
       E_reg(23) => Dangling_Input_Signal,
       E_reg(24) => Dangling_Input_Signal,
       E_reg(25) => Dangling_Input_Signal,
       E_reg(26) => Dangling_Input_Signal,
       E_reg(27) => Dangling_Input_Signal,
       E_reg(28) => Dangling_Input_Signal,
       E_reg(29) => Dangling_Input_Signal,
       E_reg(30) => Dangling_Input_Signal,
       E_reg(31) => Dangling_Input_Signal,
       E_reg(32) => Dangling_Input_Signal,
       E_reg(33) => Dangling_Input_Signal,
       E_reg(34) => Dangling_Input_Signal,
       E_reg(35) => Dangling_Input_Signal,
       E_reg(36) => Dangling_Input_Signal,
       E_reg(37) => Dangling_Input_Signal,
       E_reg(38) => Dangling_Input_Signal,
       E_reg(39) => Dangling_Input_Signal,
       E_reg(40) => Dangling_Input_Signal,
       E_reg(41) => Dangling_Input_Signal,
       E_reg(42) => Dangling_Input_Signal,
       E_reg(43) => Dangling_Input_Signal,
       E_reg(44) => Dangling_Input_Signal,
       E_reg(45) => Dangling_Input_Signal,
       E_reg(46) => Dangling_Input_Signal,
       E_reg(47) => Dangling_Input_Signal,
       E_reg(48) => Dangling_Input_Signal,
       E_reg(49) => Dangling_Input_Signal,
       E_reg(50) => Dangling_Input_Signal,
       E_reg(51) => Dangling_Input_Signal,
       E_reg(52) => Dangling_Input_Signal,
       E_reg(53) => Dangling_Input_Signal,
       E_reg(54) => Dangling_Input_Signal,
       E_reg(55) => Dangling_Input_Signal,
       E_reg(56) => Dangling_Input_Signal,
       E_reg(57) => Dangling_Input_Signal,
       E_reg(58) => Dangling_Input_Signal,
       E_reg(59) => Dangling_Input_Signal,
       E_reg(60) => Dangling_Input_Signal,
       E_reg(61) => Dangling_Input_Signal,
       E_reg(62) => Dangling_Input_Signal,
       E_reg(63) => Dangling_Input_Signal,
       E_reg(64) => Dangling_Input_Signal,
       E_reg(65) => Dangling_Input_Signal,
       E_reg(66) => Dangling_Input_Signal,
       E_reg(67) => Dangling_Input_Signal,
       E_reg(68) => Dangling_Input_Signal,
       E_reg(69) => Dangling_Input_Signal,
       E_reg(70) => Dangling_Input_Signal,
       E_reg(71) => Dangling_Input_Signal,
       E_reg(72) => Dangling_Input_Signal,
       E_reg(73) => Dangling_Input_Signal,
       E_reg(74) => Dangling_Input_Signal,
       E_reg(75) => Dangling_Input_Signal,
       E_reg(76) => Dangling_Input_Signal,
       E_reg(77) => Dangling_Input_Signal,
       E_reg(78) => Dangling_Input_Signal,
       E_reg(79) => Dangling_Input_Signal,
       E_reg(80) => Dangling_Input_Signal,
       E_reg(81) => Dangling_Input_Signal,
       E_reg(82) => Dangling_Input_Signal,
       E_reg(83) => Dangling_Input_Signal,
       E_reg(84) => Dangling_Input_Signal,
       E_reg(85) => Dangling_Input_Signal,
       E_reg(86) => Dangling_Input_Signal,
       E_reg(87) => Dangling_Input_Signal,
       E_reg(88) => Dangling_Input_Signal,
       E_reg(89) => Dangling_Input_Signal,
       E_reg(90) => Dangling_Input_Signal,
       E_reg(91) => Dangling_Input_Signal,
       E_reg(92) => Dangling_Input_Signal,
       E_reg(93) => Dangling_Input_Signal,
       E_reg(94) => Dangling_Input_Signal,
       E_reg(95) => Dangling_Input_Signal,
       E_reg(96) => Dangling_Input_Signal,
       E_reg(97) => Dangling_Input_Signal,
       E_reg(98) => Dangling_Input_Signal,
       E_reg(99) => Dangling_Input_Signal,
       E_reg(100) => Dangling_Input_Signal,
       E_reg(101) => Dangling_Input_Signal,
       E_reg(102) => Dangling_Input_Signal,
       E_reg(103) => Dangling_Input_Signal,
       E_reg(104) => Dangling_Input_Signal,
       E_reg(105) => Dangling_Input_Signal,
       E_reg(106) => Dangling_Input_Signal,
       E_reg(107) => Dangling_Input_Signal,
       E_reg(108) => Dangling_Input_Signal,
       E_reg(109) => Dangling_Input_Signal,
       E_reg(110) => Dangling_Input_Signal,
       E_reg(111) => Dangling_Input_Signal,
       E_reg(112) => Dangling_Input_Signal,
       E_reg(113) => Dangling_Input_Signal,
       E_reg(114) => Dangling_Input_Signal,
       E_reg(115) => Dangling_Input_Signal,
       E_reg(116) => Dangling_Input_Signal,
       E_reg(117) => Dangling_Input_Signal,
       E_reg(118) => Dangling_Input_Signal,
       E_reg(119) => Dangling_Input_Signal,
       E_reg(120) => Dangling_Input_Signal,
       E_reg(121) => Dangling_Input_Signal,
       E_reg(122) => Dangling_Input_Signal,
       E_reg(123) => Dangling_Input_Signal,
       E_reg(124) => Dangling_Input_Signal,
       E_reg(125) => Dangling_Input_Signal,
       E_reg(126) => Dangling_Input_Signal,
       E_reg(127) => Dangling_Input_Signal,
       F_reg(0) => Dangling_Input_Signal,
       F_reg(1) => Dangling_Input_Signal,
       F_reg(2) => Dangling_Input_Signal,
       F_reg(3) => Dangling_Input_Signal,
       F_reg(4) => Dangling_Input_Signal,
       F_reg(5) => Dangling_Input_Signal,
       F_reg(6) => Dangling_Input_Signal,
       F_reg(7) => Dangling_Input_Signal,
       F_reg(8) => Dangling_Input_Signal,
       F_reg(9) => Dangling_Input_Signal,
       F_reg(10) => Dangling_Input_Signal,
       F_reg(11) => Dangling_Input_Signal,
       F_reg(12) => Dangling_Input_Signal,
       F_reg(13) => Dangling_Input_Signal,
       F_reg(14) => Dangling_Input_Signal,
       F_reg(15) => Dangling_Input_Signal,
       F_reg(16) => Dangling_Input_Signal,
       F_reg(17) => Dangling_Input_Signal,
       F_reg(18) => Dangling_Input_Signal,
       F_reg(19) => Dangling_Input_Signal,
       F_reg(20) => Dangling_Input_Signal,
       F_reg(21) => Dangling_Input_Signal,
       F_reg(22) => Dangling_Input_Signal,
       F_reg(23) => Dangling_Input_Signal,
       F_reg(24) => Dangling_Input_Signal,
       F_reg(25) => Dangling_Input_Signal,
       F_reg(26) => Dangling_Input_Signal,
       F_reg(27) => Dangling_Input_Signal,
       F_reg(28) => Dangling_Input_Signal,
       F_reg(29) => Dangling_Input_Signal,
       F_reg(30) => Dangling_Input_Signal,
       F_reg(31) => Dangling_Input_Signal,
       F_reg(32) => Dangling_Input_Signal,
       F_reg(33) => Dangling_Input_Signal,
       F_reg(34) => Dangling_Input_Signal,
       F_reg(35) => Dangling_Input_Signal,
       F_reg(36) => Dangling_Input_Signal,
       F_reg(37) => Dangling_Input_Signal,
       F_reg(38) => Dangling_Input_Signal,
       F_reg(39) => Dangling_Input_Signal,
       F_reg(40) => Dangling_Input_Signal,
       F_reg(41) => Dangling_Input_Signal,
       F_reg(42) => Dangling_Input_Signal,
       F_reg(43) => Dangling_Input_Signal,
       F_reg(44) => Dangling_Input_Signal,
       F_reg(45) => Dangling_Input_Signal,
       F_reg(46) => Dangling_Input_Signal,
       F_reg(47) => Dangling_Input_Signal,
       F_reg(48) => Dangling_Input_Signal,
       F_reg(49) => Dangling_Input_Signal,
       F_reg(50) => Dangling_Input_Signal,
       F_reg(51) => Dangling_Input_Signal,
       F_reg(52) => Dangling_Input_Signal,
       F_reg(53) => Dangling_Input_Signal,
       F_reg(54) => Dangling_Input_Signal,
       F_reg(55) => Dangling_Input_Signal,
       F_reg(56) => Dangling_Input_Signal,
       F_reg(57) => Dangling_Input_Signal,
       F_reg(58) => Dangling_Input_Signal,
       F_reg(59) => Dangling_Input_Signal,
       F_reg(60) => Dangling_Input_Signal,
       F_reg(61) => Dangling_Input_Signal,
       F_reg(62) => Dangling_Input_Signal,
       F_reg(63) => Dangling_Input_Signal,
       F_reg(64) => Dangling_Input_Signal,
       F_reg(65) => Dangling_Input_Signal,
       F_reg(66) => Dangling_Input_Signal,
       F_reg(67) => Dangling_Input_Signal,
       F_reg(68) => Dangling_Input_Signal,
       F_reg(69) => Dangling_Input_Signal,
       F_reg(70) => Dangling_Input_Signal,
       F_reg(71) => Dangling_Input_Signal,
       F_reg(72) => Dangling_Input_Signal,
       F_reg(73) => Dangling_Input_Signal,
       F_reg(74) => Dangling_Input_Signal,
       F_reg(75) => Dangling_Input_Signal,
       F_reg(76) => Dangling_Input_Signal,
       F_reg(77) => Dangling_Input_Signal,
       F_reg(78) => Dangling_Input_Signal,
       F_reg(79) => Dangling_Input_Signal,
       F_reg(80) => Dangling_Input_Signal,
       F_reg(81) => Dangling_Input_Signal,
       F_reg(82) => Dangling_Input_Signal,
       F_reg(83) => Dangling_Input_Signal,
       F_reg(84) => Dangling_Input_Signal,
       F_reg(85) => Dangling_Input_Signal,
       F_reg(86) => Dangling_Input_Signal,
       F_reg(87) => Dangling_Input_Signal,
       F_reg(88) => Dangling_Input_Signal,
       F_reg(89) => Dangling_Input_Signal,
       F_reg(90) => Dangling_Input_Signal,
       F_reg(91) => Dangling_Input_Signal,
       F_reg(92) => Dangling_Input_Signal,
       F_reg(93) => Dangling_Input_Signal,
       F_reg(94) => Dangling_Input_Signal,
       F_reg(95) => Dangling_Input_Signal,
       F_reg(96) => Dangling_Input_Signal,
       F_reg(97) => Dangling_Input_Signal,
       F_reg(98) => Dangling_Input_Signal,
       F_reg(99) => Dangling_Input_Signal,
       F_reg(100) => Dangling_Input_Signal,
       F_reg(101) => Dangling_Input_Signal,
       F_reg(102) => Dangling_Input_Signal,
       F_reg(103) => Dangling_Input_Signal,
       F_reg(104) => Dangling_Input_Signal,
       F_reg(105) => Dangling_Input_Signal,
       F_reg(106) => Dangling_Input_Signal,
       F_reg(107) => Dangling_Input_Signal,
       F_reg(108) => Dangling_Input_Signal,
       F_reg(109) => Dangling_Input_Signal,
       F_reg(110) => Dangling_Input_Signal,
       F_reg(111) => Dangling_Input_Signal,
       F_reg(112) => Dangling_Input_Signal,
       F_reg(113) => Dangling_Input_Signal,
       F_reg(114) => Dangling_Input_Signal,
       F_reg(115) => Dangling_Input_Signal,
       F_reg(116) => Dangling_Input_Signal,
       F_reg(117) => Dangling_Input_Signal,
       F_reg(118) => Dangling_Input_Signal,
       F_reg(119) => Dangling_Input_Signal,
       F_reg(120) => Dangling_Input_Signal,
       F_reg(121) => Dangling_Input_Signal,
       F_reg(122) => Dangling_Input_Signal,
       F_reg(123) => Dangling_Input_Signal,
       F_reg(124) => Dangling_Input_Signal,
       F_reg(125) => Dangling_Input_Signal,
       F_reg(126) => Dangling_Input_Signal,
       F_reg(127) => Dangling_Input_Signal,
       odd1_Latency(0) => Dangling_Input_Signal,
       odd1_Latency(1) => Dangling_Input_Signal,
       odd1_Latency(2) => Dangling_Input_Signal,
       odd1_RegDst(0) => Dangling_Input_Signal,
       odd1_RegDst(1) => Dangling_Input_Signal,
       odd1_RegDst(2) => Dangling_Input_Signal,
       odd1_RegDst(3) => Dangling_Input_Signal,
       odd1_RegDst(4) => Dangling_Input_Signal,
       odd1_RegDst(5) => Dangling_Input_Signal,
       odd1_RegDst(6) => Dangling_Input_Signal,
       odd1_Result(0) => Dangling_Input_Signal,
       odd1_Result(1) => Dangling_Input_Signal,
       odd1_Result(2) => Dangling_Input_Signal,
       odd1_Result(3) => Dangling_Input_Signal,
       odd1_Result(4) => Dangling_Input_Signal,
       odd1_Result(5) => Dangling_Input_Signal,
       odd1_Result(6) => Dangling_Input_Signal,
       odd1_Result(7) => Dangling_Input_Signal,
       odd1_Result(8) => Dangling_Input_Signal,
       odd1_Result(9) => Dangling_Input_Signal,
       odd1_Result(10) => Dangling_Input_Signal,
       odd1_Result(11) => Dangling_Input_Signal,
       odd1_Result(12) => Dangling_Input_Signal,
       odd1_Result(13) => Dangling_Input_Signal,
       odd1_Result(14) => Dangling_Input_Signal,
       odd1_Result(15) => Dangling_Input_Signal,
       odd1_Result(16) => Dangling_Input_Signal,
       odd1_Result(17) => Dangling_Input_Signal,
       odd1_Result(18) => Dangling_Input_Signal,
       odd1_Result(19) => Dangling_Input_Signal,
       odd1_Result(20) => Dangling_Input_Signal,
       odd1_Result(21) => Dangling_Input_Signal,
       odd1_Result(22) => Dangling_Input_Signal,
       odd1_Result(23) => Dangling_Input_Signal,
       odd1_Result(24) => Dangling_Input_Signal,
       odd1_Result(25) => Dangling_Input_Signal,
       odd1_Result(26) => Dangling_Input_Signal,
       odd1_Result(27) => Dangling_Input_Signal,
       odd1_Result(28) => Dangling_Input_Signal,
       odd1_Result(29) => Dangling_Input_Signal,
       odd1_Result(30) => Dangling_Input_Signal,
       odd1_Result(31) => Dangling_Input_Signal,
       odd1_Result(32) => Dangling_Input_Signal,
       odd1_Result(33) => Dangling_Input_Signal,
       odd1_Result(34) => Dangling_Input_Signal,
       odd1_Result(35) => Dangling_Input_Signal,
       odd1_Result(36) => Dangling_Input_Signal,
       odd1_Result(37) => Dangling_Input_Signal,
       odd1_Result(38) => Dangling_Input_Signal,
       odd1_Result(39) => Dangling_Input_Signal,
       odd1_Result(40) => Dangling_Input_Signal,
       odd1_Result(41) => Dangling_Input_Signal,
       odd1_Result(42) => Dangling_Input_Signal,
       odd1_Result(43) => Dangling_Input_Signal,
       odd1_Result(44) => Dangling_Input_Signal,
       odd1_Result(45) => Dangling_Input_Signal,
       odd1_Result(46) => Dangling_Input_Signal,
       odd1_Result(47) => Dangling_Input_Signal,
       odd1_Result(48) => Dangling_Input_Signal,
       odd1_Result(49) => Dangling_Input_Signal,
       odd1_Result(50) => Dangling_Input_Signal,
       odd1_Result(51) => Dangling_Input_Signal,
       odd1_Result(52) => Dangling_Input_Signal,
       odd1_Result(53) => Dangling_Input_Signal,
       odd1_Result(54) => Dangling_Input_Signal,
       odd1_Result(55) => Dangling_Input_Signal,
       odd1_Result(56) => Dangling_Input_Signal,
       odd1_Result(57) => Dangling_Input_Signal,
       odd1_Result(58) => Dangling_Input_Signal,
       odd1_Result(59) => Dangling_Input_Signal,
       odd1_Result(60) => Dangling_Input_Signal,
       odd1_Result(61) => Dangling_Input_Signal,
       odd1_Result(62) => Dangling_Input_Signal,
       odd1_Result(63) => Dangling_Input_Signal,
       odd1_Result(64) => Dangling_Input_Signal,
       odd1_Result(65) => Dangling_Input_Signal,
       odd1_Result(66) => Dangling_Input_Signal,
       odd1_Result(67) => Dangling_Input_Signal,
       odd1_Result(68) => Dangling_Input_Signal,
       odd1_Result(69) => Dangling_Input_Signal,
       odd1_Result(70) => Dangling_Input_Signal,
       odd1_Result(71) => Dangling_Input_Signal,
       odd1_Result(72) => Dangling_Input_Signal,
       odd1_Result(73) => Dangling_Input_Signal,
       odd1_Result(74) => Dangling_Input_Signal,
       odd1_Result(75) => Dangling_Input_Signal,
       odd1_Result(76) => Dangling_Input_Signal,
       odd1_Result(77) => Dangling_Input_Signal,
       odd1_Result(78) => Dangling_Input_Signal,
       odd1_Result(79) => Dangling_Input_Signal,
       odd1_Result(80) => Dangling_Input_Signal,
       odd1_Result(81) => Dangling_Input_Signal,
       odd1_Result(82) => Dangling_Input_Signal,
       odd1_Result(83) => Dangling_Input_Signal,
       odd1_Result(84) => Dangling_Input_Signal,
       odd1_Result(85) => Dangling_Input_Signal,
       odd1_Result(86) => Dangling_Input_Signal,
       odd1_Result(87) => Dangling_Input_Signal,
       odd1_Result(88) => Dangling_Input_Signal,
       odd1_Result(89) => Dangling_Input_Signal,
       odd1_Result(90) => Dangling_Input_Signal,
       odd1_Result(91) => Dangling_Input_Signal,
       odd1_Result(92) => Dangling_Input_Signal,
       odd1_Result(93) => Dangling_Input_Signal,
       odd1_Result(94) => Dangling_Input_Signal,
       odd1_Result(95) => Dangling_Input_Signal,
       odd1_Result(96) => Dangling_Input_Signal,
       odd1_Result(97) => Dangling_Input_Signal,
       odd1_Result(98) => Dangling_Input_Signal,
       odd1_Result(99) => Dangling_Input_Signal,
       odd1_Result(100) => Dangling_Input_Signal,
       odd1_Result(101) => Dangling_Input_Signal,
       odd1_Result(102) => Dangling_Input_Signal,
       odd1_Result(103) => Dangling_Input_Signal,
       odd1_Result(104) => Dangling_Input_Signal,
       odd1_Result(105) => Dangling_Input_Signal,
       odd1_Result(106) => Dangling_Input_Signal,
       odd1_Result(107) => Dangling_Input_Signal,
       odd1_Result(108) => Dangling_Input_Signal,
       odd1_Result(109) => Dangling_Input_Signal,
       odd1_Result(110) => Dangling_Input_Signal,
       odd1_Result(111) => Dangling_Input_Signal,
       odd1_Result(112) => Dangling_Input_Signal,
       odd1_Result(113) => Dangling_Input_Signal,
       odd1_Result(114) => Dangling_Input_Signal,
       odd1_Result(115) => Dangling_Input_Signal,
       odd1_Result(116) => Dangling_Input_Signal,
       odd1_Result(117) => Dangling_Input_Signal,
       odd1_Result(118) => Dangling_Input_Signal,
       odd1_Result(119) => Dangling_Input_Signal,
       odd1_Result(120) => Dangling_Input_Signal,
       odd1_Result(121) => Dangling_Input_Signal,
       odd1_Result(122) => Dangling_Input_Signal,
       odd1_Result(123) => Dangling_Input_Signal,
       odd1_Result(124) => Dangling_Input_Signal,
       odd1_Result(125) => Dangling_Input_Signal,
       odd1_Result(126) => Dangling_Input_Signal,
       odd1_Result(127) => Dangling_Input_Signal,
       odd2_Latency(0) => Dangling_Input_Signal,
       odd2_Latency(1) => Dangling_Input_Signal,
       odd2_Latency(2) => Dangling_Input_Signal,
       odd2_RegDst(0) => Dangling_Input_Signal,
       odd2_RegDst(1) => Dangling_Input_Signal,
       odd2_RegDst(2) => Dangling_Input_Signal,
       odd2_RegDst(3) => Dangling_Input_Signal,
       odd2_RegDst(4) => Dangling_Input_Signal,
       odd2_RegDst(5) => Dangling_Input_Signal,
       odd2_RegDst(6) => Dangling_Input_Signal,
       odd2_Result(0) => Dangling_Input_Signal,
       odd2_Result(1) => Dangling_Input_Signal,
       odd2_Result(2) => Dangling_Input_Signal,
       odd2_Result(3) => Dangling_Input_Signal,
       odd2_Result(4) => Dangling_Input_Signal,
       odd2_Result(5) => Dangling_Input_Signal,
       odd2_Result(6) => Dangling_Input_Signal,
       odd2_Result(7) => Dangling_Input_Signal,
       odd2_Result(8) => Dangling_Input_Signal,
       odd2_Result(9) => Dangling_Input_Signal,
       odd2_Result(10) => Dangling_Input_Signal,
       odd2_Result(11) => Dangling_Input_Signal,
       odd2_Result(12) => Dangling_Input_Signal,
       odd2_Result(13) => Dangling_Input_Signal,
       odd2_Result(14) => Dangling_Input_Signal,
       odd2_Result(15) => Dangling_Input_Signal,
       odd2_Result(16) => Dangling_Input_Signal,
       odd2_Result(17) => Dangling_Input_Signal,
       odd2_Result(18) => Dangling_Input_Signal,
       odd2_Result(19) => Dangling_Input_Signal,
       odd2_Result(20) => Dangling_Input_Signal,
       odd2_Result(21) => Dangling_Input_Signal,
       odd2_Result(22) => Dangling_Input_Signal,
       odd2_Result(23) => Dangling_Input_Signal,
       odd2_Result(24) => Dangling_Input_Signal,
       odd2_Result(25) => Dangling_Input_Signal,
       odd2_Result(26) => Dangling_Input_Signal,
       odd2_Result(27) => Dangling_Input_Signal,
       odd2_Result(28) => Dangling_Input_Signal,
       odd2_Result(29) => Dangling_Input_Signal,
       odd2_Result(30) => Dangling_Input_Signal,
       odd2_Result(31) => Dangling_Input_Signal,
       odd2_Result(32) => Dangling_Input_Signal,
       odd2_Result(33) => Dangling_Input_Signal,
       odd2_Result(34) => Dangling_Input_Signal,
       odd2_Result(35) => Dangling_Input_Signal,
       odd2_Result(36) => Dangling_Input_Signal,
       odd2_Result(37) => Dangling_Input_Signal,
       odd2_Result(38) => Dangling_Input_Signal,
       odd2_Result(39) => Dangling_Input_Signal,
       odd2_Result(40) => Dangling_Input_Signal,
       odd2_Result(41) => Dangling_Input_Signal,
       odd2_Result(42) => Dangling_Input_Signal,
       odd2_Result(43) => Dangling_Input_Signal,
       odd2_Result(44) => Dangling_Input_Signal,
       odd2_Result(45) => Dangling_Input_Signal,
       odd2_Result(46) => Dangling_Input_Signal,
       odd2_Result(47) => Dangling_Input_Signal,
       odd2_Result(48) => Dangling_Input_Signal,
       odd2_Result(49) => Dangling_Input_Signal,
       odd2_Result(50) => Dangling_Input_Signal,
       odd2_Result(51) => Dangling_Input_Signal,
       odd2_Result(52) => Dangling_Input_Signal,
       odd2_Result(53) => Dangling_Input_Signal,
       odd2_Result(54) => Dangling_Input_Signal,
       odd2_Result(55) => Dangling_Input_Signal,
       odd2_Result(56) => Dangling_Input_Signal,
       odd2_Result(57) => Dangling_Input_Signal,
       odd2_Result(58) => Dangling_Input_Signal,
       odd2_Result(59) => Dangling_Input_Signal,
       odd2_Result(60) => Dangling_Input_Signal,
       odd2_Result(61) => Dangling_Input_Signal,
       odd2_Result(62) => Dangling_Input_Signal,
       odd2_Result(63) => Dangling_Input_Signal,
       odd2_Result(64) => Dangling_Input_Signal,
       odd2_Result(65) => Dangling_Input_Signal,
       odd2_Result(66) => Dangling_Input_Signal,
       odd2_Result(67) => Dangling_Input_Signal,
       odd2_Result(68) => Dangling_Input_Signal,
       odd2_Result(69) => Dangling_Input_Signal,
       odd2_Result(70) => Dangling_Input_Signal,
       odd2_Result(71) => Dangling_Input_Signal,
       odd2_Result(72) => Dangling_Input_Signal,
       odd2_Result(73) => Dangling_Input_Signal,
       odd2_Result(74) => Dangling_Input_Signal,
       odd2_Result(75) => Dangling_Input_Signal,
       odd2_Result(76) => Dangling_Input_Signal,
       odd2_Result(77) => Dangling_Input_Signal,
       odd2_Result(78) => Dangling_Input_Signal,
       odd2_Result(79) => Dangling_Input_Signal,
       odd2_Result(80) => Dangling_Input_Signal,
       odd2_Result(81) => Dangling_Input_Signal,
       odd2_Result(82) => Dangling_Input_Signal,
       odd2_Result(83) => Dangling_Input_Signal,
       odd2_Result(84) => Dangling_Input_Signal,
       odd2_Result(85) => Dangling_Input_Signal,
       odd2_Result(86) => Dangling_Input_Signal,
       odd2_Result(87) => Dangling_Input_Signal,
       odd2_Result(88) => Dangling_Input_Signal,
       odd2_Result(89) => Dangling_Input_Signal,
       odd2_Result(90) => Dangling_Input_Signal,
       odd2_Result(91) => Dangling_Input_Signal,
       odd2_Result(92) => Dangling_Input_Signal,
       odd2_Result(93) => Dangling_Input_Signal,
       odd2_Result(94) => Dangling_Input_Signal,
       odd2_Result(95) => Dangling_Input_Signal,
       odd2_Result(96) => Dangling_Input_Signal,
       odd2_Result(97) => Dangling_Input_Signal,
       odd2_Result(98) => Dangling_Input_Signal,
       odd2_Result(99) => Dangling_Input_Signal,
       odd2_Result(100) => Dangling_Input_Signal,
       odd2_Result(101) => Dangling_Input_Signal,
       odd2_Result(102) => Dangling_Input_Signal,
       odd2_Result(103) => Dangling_Input_Signal,
       odd2_Result(104) => Dangling_Input_Signal,
       odd2_Result(105) => Dangling_Input_Signal,
       odd2_Result(106) => Dangling_Input_Signal,
       odd2_Result(107) => Dangling_Input_Signal,
       odd2_Result(108) => Dangling_Input_Signal,
       odd2_Result(109) => Dangling_Input_Signal,
       odd2_Result(110) => Dangling_Input_Signal,
       odd2_Result(111) => Dangling_Input_Signal,
       odd2_Result(112) => Dangling_Input_Signal,
       odd2_Result(113) => Dangling_Input_Signal,
       odd2_Result(114) => Dangling_Input_Signal,
       odd2_Result(115) => Dangling_Input_Signal,
       odd2_Result(116) => Dangling_Input_Signal,
       odd2_Result(117) => Dangling_Input_Signal,
       odd2_Result(118) => Dangling_Input_Signal,
       odd2_Result(119) => Dangling_Input_Signal,
       odd2_Result(120) => Dangling_Input_Signal,
       odd2_Result(121) => Dangling_Input_Signal,
       odd2_Result(122) => Dangling_Input_Signal,
       odd2_Result(123) => Dangling_Input_Signal,
       odd2_Result(124) => Dangling_Input_Signal,
       odd2_Result(125) => Dangling_Input_Signal,
       odd2_Result(126) => Dangling_Input_Signal,
       odd2_Result(127) => Dangling_Input_Signal,
       odd3_Latency(0) => Dangling_Input_Signal,
       odd3_Latency(1) => Dangling_Input_Signal,
       odd3_Latency(2) => Dangling_Input_Signal,
       odd3_RegDst(0) => Dangling_Input_Signal,
       odd3_RegDst(1) => Dangling_Input_Signal,
       odd3_RegDst(2) => Dangling_Input_Signal,
       odd3_RegDst(3) => Dangling_Input_Signal,
       odd3_RegDst(4) => Dangling_Input_Signal,
       odd3_RegDst(5) => Dangling_Input_Signal,
       odd3_RegDst(6) => Dangling_Input_Signal,
       odd3_Result(0) => Dangling_Input_Signal,
       odd3_Result(1) => Dangling_Input_Signal,
       odd3_Result(2) => Dangling_Input_Signal,
       odd3_Result(3) => Dangling_Input_Signal,
       odd3_Result(4) => Dangling_Input_Signal,
       odd3_Result(5) => Dangling_Input_Signal,
       odd3_Result(6) => Dangling_Input_Signal,
       odd3_Result(7) => Dangling_Input_Signal,
       odd3_Result(8) => Dangling_Input_Signal,
       odd3_Result(9) => Dangling_Input_Signal,
       odd3_Result(10) => Dangling_Input_Signal,
       odd3_Result(11) => Dangling_Input_Signal,
       odd3_Result(12) => Dangling_Input_Signal,
       odd3_Result(13) => Dangling_Input_Signal,
       odd3_Result(14) => Dangling_Input_Signal,
       odd3_Result(15) => Dangling_Input_Signal,
       odd3_Result(16) => Dangling_Input_Signal,
       odd3_Result(17) => Dangling_Input_Signal,
       odd3_Result(18) => Dangling_Input_Signal,
       odd3_Result(19) => Dangling_Input_Signal,
       odd3_Result(20) => Dangling_Input_Signal,
       odd3_Result(21) => Dangling_Input_Signal,
       odd3_Result(22) => Dangling_Input_Signal,
       odd3_Result(23) => Dangling_Input_Signal,
       odd3_Result(24) => Dangling_Input_Signal,
       odd3_Result(25) => Dangling_Input_Signal,
       odd3_Result(26) => Dangling_Input_Signal,
       odd3_Result(27) => Dangling_Input_Signal,
       odd3_Result(28) => Dangling_Input_Signal,
       odd3_Result(29) => Dangling_Input_Signal,
       odd3_Result(30) => Dangling_Input_Signal,
       odd3_Result(31) => Dangling_Input_Signal,
       odd3_Result(32) => Dangling_Input_Signal,
       odd3_Result(33) => Dangling_Input_Signal,
       odd3_Result(34) => Dangling_Input_Signal,
       odd3_Result(35) => Dangling_Input_Signal,
       odd3_Result(36) => Dangling_Input_Signal,
       odd3_Result(37) => Dangling_Input_Signal,
       odd3_Result(38) => Dangling_Input_Signal,
       odd3_Result(39) => Dangling_Input_Signal,
       odd3_Result(40) => Dangling_Input_Signal,
       odd3_Result(41) => Dangling_Input_Signal,
       odd3_Result(42) => Dangling_Input_Signal,
       odd3_Result(43) => Dangling_Input_Signal,
       odd3_Result(44) => Dangling_Input_Signal,
       odd3_Result(45) => Dangling_Input_Signal,
       odd3_Result(46) => Dangling_Input_Signal,
       odd3_Result(47) => Dangling_Input_Signal,
       odd3_Result(48) => Dangling_Input_Signal,
       odd3_Result(49) => Dangling_Input_Signal,
       odd3_Result(50) => Dangling_Input_Signal,
       odd3_Result(51) => Dangling_Input_Signal,
       odd3_Result(52) => Dangling_Input_Signal,
       odd3_Result(53) => Dangling_Input_Signal,
       odd3_Result(54) => Dangling_Input_Signal,
       odd3_Result(55) => Dangling_Input_Signal,
       odd3_Result(56) => Dangling_Input_Signal,
       odd3_Result(57) => Dangling_Input_Signal,
       odd3_Result(58) => Dangling_Input_Signal,
       odd3_Result(59) => Dangling_Input_Signal,
       odd3_Result(60) => Dangling_Input_Signal,
       odd3_Result(61) => Dangling_Input_Signal,
       odd3_Result(62) => Dangling_Input_Signal,
       odd3_Result(63) => Dangling_Input_Signal,
       odd3_Result(64) => Dangling_Input_Signal,
       odd3_Result(65) => Dangling_Input_Signal,
       odd3_Result(66) => Dangling_Input_Signal,
       odd3_Result(67) => Dangling_Input_Signal,
       odd3_Result(68) => Dangling_Input_Signal,
       odd3_Result(69) => Dangling_Input_Signal,
       odd3_Result(70) => Dangling_Input_Signal,
       odd3_Result(71) => Dangling_Input_Signal,
       odd3_Result(72) => Dangling_Input_Signal,
       odd3_Result(73) => Dangling_Input_Signal,
       odd3_Result(74) => Dangling_Input_Signal,
       odd3_Result(75) => Dangling_Input_Signal,
       odd3_Result(76) => Dangling_Input_Signal,
       odd3_Result(77) => Dangling_Input_Signal,
       odd3_Result(78) => Dangling_Input_Signal,
       odd3_Result(79) => Dangling_Input_Signal,
       odd3_Result(80) => Dangling_Input_Signal,
       odd3_Result(81) => Dangling_Input_Signal,
       odd3_Result(82) => Dangling_Input_Signal,
       odd3_Result(83) => Dangling_Input_Signal,
       odd3_Result(84) => Dangling_Input_Signal,
       odd3_Result(85) => Dangling_Input_Signal,
       odd3_Result(86) => Dangling_Input_Signal,
       odd3_Result(87) => Dangling_Input_Signal,
       odd3_Result(88) => Dangling_Input_Signal,
       odd3_Result(89) => Dangling_Input_Signal,
       odd3_Result(90) => Dangling_Input_Signal,
       odd3_Result(91) => Dangling_Input_Signal,
       odd3_Result(92) => Dangling_Input_Signal,
       odd3_Result(93) => Dangling_Input_Signal,
       odd3_Result(94) => Dangling_Input_Signal,
       odd3_Result(95) => Dangling_Input_Signal,
       odd3_Result(96) => Dangling_Input_Signal,
       odd3_Result(97) => Dangling_Input_Signal,
       odd3_Result(98) => Dangling_Input_Signal,
       odd3_Result(99) => Dangling_Input_Signal,
       odd3_Result(100) => Dangling_Input_Signal,
       odd3_Result(101) => Dangling_Input_Signal,
       odd3_Result(102) => Dangling_Input_Signal,
       odd3_Result(103) => Dangling_Input_Signal,
       odd3_Result(104) => Dangling_Input_Signal,
       odd3_Result(105) => Dangling_Input_Signal,
       odd3_Result(106) => Dangling_Input_Signal,
       odd3_Result(107) => Dangling_Input_Signal,
       odd3_Result(108) => Dangling_Input_Signal,
       odd3_Result(109) => Dangling_Input_Signal,
       odd3_Result(110) => Dangling_Input_Signal,
       odd3_Result(111) => Dangling_Input_Signal,
       odd3_Result(112) => Dangling_Input_Signal,
       odd3_Result(113) => Dangling_Input_Signal,
       odd3_Result(114) => Dangling_Input_Signal,
       odd3_Result(115) => Dangling_Input_Signal,
       odd3_Result(116) => Dangling_Input_Signal,
       odd3_Result(117) => Dangling_Input_Signal,
       odd3_Result(118) => Dangling_Input_Signal,
       odd3_Result(119) => Dangling_Input_Signal,
       odd3_Result(120) => Dangling_Input_Signal,
       odd3_Result(121) => Dangling_Input_Signal,
       odd3_Result(122) => Dangling_Input_Signal,
       odd3_Result(123) => Dangling_Input_Signal,
       odd3_Result(124) => Dangling_Input_Signal,
       odd3_Result(125) => Dangling_Input_Signal,
       odd3_Result(126) => Dangling_Input_Signal,
       odd3_Result(127) => Dangling_Input_Signal,
       odd4_Latency(0) => Dangling_Input_Signal,
       odd4_Latency(1) => Dangling_Input_Signal,
       odd4_Latency(2) => Dangling_Input_Signal,
       odd4_RegDst(0) => Dangling_Input_Signal,
       odd4_RegDst(1) => Dangling_Input_Signal,
       odd4_RegDst(2) => Dangling_Input_Signal,
       odd4_RegDst(3) => Dangling_Input_Signal,
       odd4_RegDst(4) => Dangling_Input_Signal,
       odd4_RegDst(5) => Dangling_Input_Signal,
       odd4_RegDst(6) => Dangling_Input_Signal,
       odd4_Result(0) => Dangling_Input_Signal,
       odd4_Result(1) => Dangling_Input_Signal,
       odd4_Result(2) => Dangling_Input_Signal,
       odd4_Result(3) => Dangling_Input_Signal,
       odd4_Result(4) => Dangling_Input_Signal,
       odd4_Result(5) => Dangling_Input_Signal,
       odd4_Result(6) => Dangling_Input_Signal,
       odd4_Result(7) => Dangling_Input_Signal,
       odd4_Result(8) => Dangling_Input_Signal,
       odd4_Result(9) => Dangling_Input_Signal,
       odd4_Result(10) => Dangling_Input_Signal,
       odd4_Result(11) => Dangling_Input_Signal,
       odd4_Result(12) => Dangling_Input_Signal,
       odd4_Result(13) => Dangling_Input_Signal,
       odd4_Result(14) => Dangling_Input_Signal,
       odd4_Result(15) => Dangling_Input_Signal,
       odd4_Result(16) => Dangling_Input_Signal,
       odd4_Result(17) => Dangling_Input_Signal,
       odd4_Result(18) => Dangling_Input_Signal,
       odd4_Result(19) => Dangling_Input_Signal,
       odd4_Result(20) => Dangling_Input_Signal,
       odd4_Result(21) => Dangling_Input_Signal,
       odd4_Result(22) => Dangling_Input_Signal,
       odd4_Result(23) => Dangling_Input_Signal,
       odd4_Result(24) => Dangling_Input_Signal,
       odd4_Result(25) => Dangling_Input_Signal,
       odd4_Result(26) => Dangling_Input_Signal,
       odd4_Result(27) => Dangling_Input_Signal,
       odd4_Result(28) => Dangling_Input_Signal,
       odd4_Result(29) => Dangling_Input_Signal,
       odd4_Result(30) => Dangling_Input_Signal,
       odd4_Result(31) => Dangling_Input_Signal,
       odd4_Result(32) => Dangling_Input_Signal,
       odd4_Result(33) => Dangling_Input_Signal,
       odd4_Result(34) => Dangling_Input_Signal,
       odd4_Result(35) => Dangling_Input_Signal,
       odd4_Result(36) => Dangling_Input_Signal,
       odd4_Result(37) => Dangling_Input_Signal,
       odd4_Result(38) => Dangling_Input_Signal,
       odd4_Result(39) => Dangling_Input_Signal,
       odd4_Result(40) => Dangling_Input_Signal,
       odd4_Result(41) => Dangling_Input_Signal,
       odd4_Result(42) => Dangling_Input_Signal,
       odd4_Result(43) => Dangling_Input_Signal,
       odd4_Result(44) => Dangling_Input_Signal,
       odd4_Result(45) => Dangling_Input_Signal,
       odd4_Result(46) => Dangling_Input_Signal,
       odd4_Result(47) => Dangling_Input_Signal,
       odd4_Result(48) => Dangling_Input_Signal,
       odd4_Result(49) => Dangling_Input_Signal,
       odd4_Result(50) => Dangling_Input_Signal,
       odd4_Result(51) => Dangling_Input_Signal,
       odd4_Result(52) => Dangling_Input_Signal,
       odd4_Result(53) => Dangling_Input_Signal,
       odd4_Result(54) => Dangling_Input_Signal,
       odd4_Result(55) => Dangling_Input_Signal,
       odd4_Result(56) => Dangling_Input_Signal,
       odd4_Result(57) => Dangling_Input_Signal,
       odd4_Result(58) => Dangling_Input_Signal,
       odd4_Result(59) => Dangling_Input_Signal,
       odd4_Result(60) => Dangling_Input_Signal,
       odd4_Result(61) => Dangling_Input_Signal,
       odd4_Result(62) => Dangling_Input_Signal,
       odd4_Result(63) => Dangling_Input_Signal,
       odd4_Result(64) => Dangling_Input_Signal,
       odd4_Result(65) => Dangling_Input_Signal,
       odd4_Result(66) => Dangling_Input_Signal,
       odd4_Result(67) => Dangling_Input_Signal,
       odd4_Result(68) => Dangling_Input_Signal,
       odd4_Result(69) => Dangling_Input_Signal,
       odd4_Result(70) => Dangling_Input_Signal,
       odd4_Result(71) => Dangling_Input_Signal,
       odd4_Result(72) => Dangling_Input_Signal,
       odd4_Result(73) => Dangling_Input_Signal,
       odd4_Result(74) => Dangling_Input_Signal,
       odd4_Result(75) => Dangling_Input_Signal,
       odd4_Result(76) => Dangling_Input_Signal,
       odd4_Result(77) => Dangling_Input_Signal,
       odd4_Result(78) => Dangling_Input_Signal,
       odd4_Result(79) => Dangling_Input_Signal,
       odd4_Result(80) => Dangling_Input_Signal,
       odd4_Result(81) => Dangling_Input_Signal,
       odd4_Result(82) => Dangling_Input_Signal,
       odd4_Result(83) => Dangling_Input_Signal,
       odd4_Result(84) => Dangling_Input_Signal,
       odd4_Result(85) => Dangling_Input_Signal,
       odd4_Result(86) => Dangling_Input_Signal,
       odd4_Result(87) => Dangling_Input_Signal,
       odd4_Result(88) => Dangling_Input_Signal,
       odd4_Result(89) => Dangling_Input_Signal,
       odd4_Result(90) => Dangling_Input_Signal,
       odd4_Result(91) => Dangling_Input_Signal,
       odd4_Result(92) => Dangling_Input_Signal,
       odd4_Result(93) => Dangling_Input_Signal,
       odd4_Result(94) => Dangling_Input_Signal,
       odd4_Result(95) => Dangling_Input_Signal,
       odd4_Result(96) => Dangling_Input_Signal,
       odd4_Result(97) => Dangling_Input_Signal,
       odd4_Result(98) => Dangling_Input_Signal,
       odd4_Result(99) => Dangling_Input_Signal,
       odd4_Result(100) => Dangling_Input_Signal,
       odd4_Result(101) => Dangling_Input_Signal,
       odd4_Result(102) => Dangling_Input_Signal,
       odd4_Result(103) => Dangling_Input_Signal,
       odd4_Result(104) => Dangling_Input_Signal,
       odd4_Result(105) => Dangling_Input_Signal,
       odd4_Result(106) => Dangling_Input_Signal,
       odd4_Result(107) => Dangling_Input_Signal,
       odd4_Result(108) => Dangling_Input_Signal,
       odd4_Result(109) => Dangling_Input_Signal,
       odd4_Result(110) => Dangling_Input_Signal,
       odd4_Result(111) => Dangling_Input_Signal,
       odd4_Result(112) => Dangling_Input_Signal,
       odd4_Result(113) => Dangling_Input_Signal,
       odd4_Result(114) => Dangling_Input_Signal,
       odd4_Result(115) => Dangling_Input_Signal,
       odd4_Result(116) => Dangling_Input_Signal,
       odd4_Result(117) => Dangling_Input_Signal,
       odd4_Result(118) => Dangling_Input_Signal,
       odd4_Result(119) => Dangling_Input_Signal,
       odd4_Result(120) => Dangling_Input_Signal,
       odd4_Result(121) => Dangling_Input_Signal,
       odd4_Result(122) => Dangling_Input_Signal,
       odd4_Result(123) => Dangling_Input_Signal,
       odd4_Result(124) => Dangling_Input_Signal,
       odd4_Result(125) => Dangling_Input_Signal,
       odd4_Result(126) => Dangling_Input_Signal,
       odd4_Result(127) => Dangling_Input_Signal,
       odd5_Latency(0) => Dangling_Input_Signal,
       odd5_Latency(1) => Dangling_Input_Signal,
       odd5_Latency(2) => Dangling_Input_Signal,
       odd5_RegDst(0) => Dangling_Input_Signal,
       odd5_RegDst(1) => Dangling_Input_Signal,
       odd5_RegDst(2) => Dangling_Input_Signal,
       odd5_RegDst(3) => Dangling_Input_Signal,
       odd5_RegDst(4) => Dangling_Input_Signal,
       odd5_RegDst(5) => Dangling_Input_Signal,
       odd5_RegDst(6) => Dangling_Input_Signal,
       odd5_Result(0) => Dangling_Input_Signal,
       odd5_Result(1) => Dangling_Input_Signal,
       odd5_Result(2) => Dangling_Input_Signal,
       odd5_Result(3) => Dangling_Input_Signal,
       odd5_Result(4) => Dangling_Input_Signal,
       odd5_Result(5) => Dangling_Input_Signal,
       odd5_Result(6) => Dangling_Input_Signal,
       odd5_Result(7) => Dangling_Input_Signal,
       odd5_Result(8) => Dangling_Input_Signal,
       odd5_Result(9) => Dangling_Input_Signal,
       odd5_Result(10) => Dangling_Input_Signal,
       odd5_Result(11) => Dangling_Input_Signal,
       odd5_Result(12) => Dangling_Input_Signal,
       odd5_Result(13) => Dangling_Input_Signal,
       odd5_Result(14) => Dangling_Input_Signal,
       odd5_Result(15) => Dangling_Input_Signal,
       odd5_Result(16) => Dangling_Input_Signal,
       odd5_Result(17) => Dangling_Input_Signal,
       odd5_Result(18) => Dangling_Input_Signal,
       odd5_Result(19) => Dangling_Input_Signal,
       odd5_Result(20) => Dangling_Input_Signal,
       odd5_Result(21) => Dangling_Input_Signal,
       odd5_Result(22) => Dangling_Input_Signal,
       odd5_Result(23) => Dangling_Input_Signal,
       odd5_Result(24) => Dangling_Input_Signal,
       odd5_Result(25) => Dangling_Input_Signal,
       odd5_Result(26) => Dangling_Input_Signal,
       odd5_Result(27) => Dangling_Input_Signal,
       odd5_Result(28) => Dangling_Input_Signal,
       odd5_Result(29) => Dangling_Input_Signal,
       odd5_Result(30) => Dangling_Input_Signal,
       odd5_Result(31) => Dangling_Input_Signal,
       odd5_Result(32) => Dangling_Input_Signal,
       odd5_Result(33) => Dangling_Input_Signal,
       odd5_Result(34) => Dangling_Input_Signal,
       odd5_Result(35) => Dangling_Input_Signal,
       odd5_Result(36) => Dangling_Input_Signal,
       odd5_Result(37) => Dangling_Input_Signal,
       odd5_Result(38) => Dangling_Input_Signal,
       odd5_Result(39) => Dangling_Input_Signal,
       odd5_Result(40) => Dangling_Input_Signal,
       odd5_Result(41) => Dangling_Input_Signal,
       odd5_Result(42) => Dangling_Input_Signal,
       odd5_Result(43) => Dangling_Input_Signal,
       odd5_Result(44) => Dangling_Input_Signal,
       odd5_Result(45) => Dangling_Input_Signal,
       odd5_Result(46) => Dangling_Input_Signal,
       odd5_Result(47) => Dangling_Input_Signal,
       odd5_Result(48) => Dangling_Input_Signal,
       odd5_Result(49) => Dangling_Input_Signal,
       odd5_Result(50) => Dangling_Input_Signal,
       odd5_Result(51) => Dangling_Input_Signal,
       odd5_Result(52) => Dangling_Input_Signal,
       odd5_Result(53) => Dangling_Input_Signal,
       odd5_Result(54) => Dangling_Input_Signal,
       odd5_Result(55) => Dangling_Input_Signal,
       odd5_Result(56) => Dangling_Input_Signal,
       odd5_Result(57) => Dangling_Input_Signal,
       odd5_Result(58) => Dangling_Input_Signal,
       odd5_Result(59) => Dangling_Input_Signal,
       odd5_Result(60) => Dangling_Input_Signal,
       odd5_Result(61) => Dangling_Input_Signal,
       odd5_Result(62) => Dangling_Input_Signal,
       odd5_Result(63) => Dangling_Input_Signal,
       odd5_Result(64) => Dangling_Input_Signal,
       odd5_Result(65) => Dangling_Input_Signal,
       odd5_Result(66) => Dangling_Input_Signal,
       odd5_Result(67) => Dangling_Input_Signal,
       odd5_Result(68) => Dangling_Input_Signal,
       odd5_Result(69) => Dangling_Input_Signal,
       odd5_Result(70) => Dangling_Input_Signal,
       odd5_Result(71) => Dangling_Input_Signal,
       odd5_Result(72) => Dangling_Input_Signal,
       odd5_Result(73) => Dangling_Input_Signal,
       odd5_Result(74) => Dangling_Input_Signal,
       odd5_Result(75) => Dangling_Input_Signal,
       odd5_Result(76) => Dangling_Input_Signal,
       odd5_Result(77) => Dangling_Input_Signal,
       odd5_Result(78) => Dangling_Input_Signal,
       odd5_Result(79) => Dangling_Input_Signal,
       odd5_Result(80) => Dangling_Input_Signal,
       odd5_Result(81) => Dangling_Input_Signal,
       odd5_Result(82) => Dangling_Input_Signal,
       odd5_Result(83) => Dangling_Input_Signal,
       odd5_Result(84) => Dangling_Input_Signal,
       odd5_Result(85) => Dangling_Input_Signal,
       odd5_Result(86) => Dangling_Input_Signal,
       odd5_Result(87) => Dangling_Input_Signal,
       odd5_Result(88) => Dangling_Input_Signal,
       odd5_Result(89) => Dangling_Input_Signal,
       odd5_Result(90) => Dangling_Input_Signal,
       odd5_Result(91) => Dangling_Input_Signal,
       odd5_Result(92) => Dangling_Input_Signal,
       odd5_Result(93) => Dangling_Input_Signal,
       odd5_Result(94) => Dangling_Input_Signal,
       odd5_Result(95) => Dangling_Input_Signal,
       odd5_Result(96) => Dangling_Input_Signal,
       odd5_Result(97) => Dangling_Input_Signal,
       odd5_Result(98) => Dangling_Input_Signal,
       odd5_Result(99) => Dangling_Input_Signal,
       odd5_Result(100) => Dangling_Input_Signal,
       odd5_Result(101) => Dangling_Input_Signal,
       odd5_Result(102) => Dangling_Input_Signal,
       odd5_Result(103) => Dangling_Input_Signal,
       odd5_Result(104) => Dangling_Input_Signal,
       odd5_Result(105) => Dangling_Input_Signal,
       odd5_Result(106) => Dangling_Input_Signal,
       odd5_Result(107) => Dangling_Input_Signal,
       odd5_Result(108) => Dangling_Input_Signal,
       odd5_Result(109) => Dangling_Input_Signal,
       odd5_Result(110) => Dangling_Input_Signal,
       odd5_Result(111) => Dangling_Input_Signal,
       odd5_Result(112) => Dangling_Input_Signal,
       odd5_Result(113) => Dangling_Input_Signal,
       odd5_Result(114) => Dangling_Input_Signal,
       odd5_Result(115) => Dangling_Input_Signal,
       odd5_Result(116) => Dangling_Input_Signal,
       odd5_Result(117) => Dangling_Input_Signal,
       odd5_Result(118) => Dangling_Input_Signal,
       odd5_Result(119) => Dangling_Input_Signal,
       odd5_Result(120) => Dangling_Input_Signal,
       odd5_Result(121) => Dangling_Input_Signal,
       odd5_Result(122) => Dangling_Input_Signal,
       odd5_Result(123) => Dangling_Input_Signal,
       odd5_Result(124) => Dangling_Input_Signal,
       odd5_Result(125) => Dangling_Input_Signal,
       odd5_Result(126) => Dangling_Input_Signal,
       odd5_Result(127) => Dangling_Input_Signal,
       odd6_Latency(0) => Dangling_Input_Signal,
       odd6_Latency(1) => Dangling_Input_Signal,
       odd6_Latency(2) => Dangling_Input_Signal,
       odd6_RegDst(0) => Dangling_Input_Signal,
       odd6_RegDst(1) => Dangling_Input_Signal,
       odd6_RegDst(2) => Dangling_Input_Signal,
       odd6_RegDst(3) => Dangling_Input_Signal,
       odd6_RegDst(4) => Dangling_Input_Signal,
       odd6_RegDst(5) => Dangling_Input_Signal,
       odd6_RegDst(6) => Dangling_Input_Signal,
       odd6_Result(0) => Dangling_Input_Signal,
       odd6_Result(1) => Dangling_Input_Signal,
       odd6_Result(2) => Dangling_Input_Signal,
       odd6_Result(3) => Dangling_Input_Signal,
       odd6_Result(4) => Dangling_Input_Signal,
       odd6_Result(5) => Dangling_Input_Signal,
       odd6_Result(6) => Dangling_Input_Signal,
       odd6_Result(7) => Dangling_Input_Signal,
       odd6_Result(8) => Dangling_Input_Signal,
       odd6_Result(9) => Dangling_Input_Signal,
       odd6_Result(10) => Dangling_Input_Signal,
       odd6_Result(11) => Dangling_Input_Signal,
       odd6_Result(12) => Dangling_Input_Signal,
       odd6_Result(13) => Dangling_Input_Signal,
       odd6_Result(14) => Dangling_Input_Signal,
       odd6_Result(15) => Dangling_Input_Signal,
       odd6_Result(16) => Dangling_Input_Signal,
       odd6_Result(17) => Dangling_Input_Signal,
       odd6_Result(18) => Dangling_Input_Signal,
       odd6_Result(19) => Dangling_Input_Signal,
       odd6_Result(20) => Dangling_Input_Signal,
       odd6_Result(21) => Dangling_Input_Signal,
       odd6_Result(22) => Dangling_Input_Signal,
       odd6_Result(23) => Dangling_Input_Signal,
       odd6_Result(24) => Dangling_Input_Signal,
       odd6_Result(25) => Dangling_Input_Signal,
       odd6_Result(26) => Dangling_Input_Signal,
       odd6_Result(27) => Dangling_Input_Signal,
       odd6_Result(28) => Dangling_Input_Signal,
       odd6_Result(29) => Dangling_Input_Signal,
       odd6_Result(30) => Dangling_Input_Signal,
       odd6_Result(31) => Dangling_Input_Signal,
       odd6_Result(32) => Dangling_Input_Signal,
       odd6_Result(33) => Dangling_Input_Signal,
       odd6_Result(34) => Dangling_Input_Signal,
       odd6_Result(35) => Dangling_Input_Signal,
       odd6_Result(36) => Dangling_Input_Signal,
       odd6_Result(37) => Dangling_Input_Signal,
       odd6_Result(38) => Dangling_Input_Signal,
       odd6_Result(39) => Dangling_Input_Signal,
       odd6_Result(40) => Dangling_Input_Signal,
       odd6_Result(41) => Dangling_Input_Signal,
       odd6_Result(42) => Dangling_Input_Signal,
       odd6_Result(43) => Dangling_Input_Signal,
       odd6_Result(44) => Dangling_Input_Signal,
       odd6_Result(45) => Dangling_Input_Signal,
       odd6_Result(46) => Dangling_Input_Signal,
       odd6_Result(47) => Dangling_Input_Signal,
       odd6_Result(48) => Dangling_Input_Signal,
       odd6_Result(49) => Dangling_Input_Signal,
       odd6_Result(50) => Dangling_Input_Signal,
       odd6_Result(51) => Dangling_Input_Signal,
       odd6_Result(52) => Dangling_Input_Signal,
       odd6_Result(53) => Dangling_Input_Signal,
       odd6_Result(54) => Dangling_Input_Signal,
       odd6_Result(55) => Dangling_Input_Signal,
       odd6_Result(56) => Dangling_Input_Signal,
       odd6_Result(57) => Dangling_Input_Signal,
       odd6_Result(58) => Dangling_Input_Signal,
       odd6_Result(59) => Dangling_Input_Signal,
       odd6_Result(60) => Dangling_Input_Signal,
       odd6_Result(61) => Dangling_Input_Signal,
       odd6_Result(62) => Dangling_Input_Signal,
       odd6_Result(63) => Dangling_Input_Signal,
       odd6_Result(64) => Dangling_Input_Signal,
       odd6_Result(65) => Dangling_Input_Signal,
       odd6_Result(66) => Dangling_Input_Signal,
       odd6_Result(67) => Dangling_Input_Signal,
       odd6_Result(68) => Dangling_Input_Signal,
       odd6_Result(69) => Dangling_Input_Signal,
       odd6_Result(70) => Dangling_Input_Signal,
       odd6_Result(71) => Dangling_Input_Signal,
       odd6_Result(72) => Dangling_Input_Signal,
       odd6_Result(73) => Dangling_Input_Signal,
       odd6_Result(74) => Dangling_Input_Signal,
       odd6_Result(75) => Dangling_Input_Signal,
       odd6_Result(76) => Dangling_Input_Signal,
       odd6_Result(77) => Dangling_Input_Signal,
       odd6_Result(78) => Dangling_Input_Signal,
       odd6_Result(79) => Dangling_Input_Signal,
       odd6_Result(80) => Dangling_Input_Signal,
       odd6_Result(81) => Dangling_Input_Signal,
       odd6_Result(82) => Dangling_Input_Signal,
       odd6_Result(83) => Dangling_Input_Signal,
       odd6_Result(84) => Dangling_Input_Signal,
       odd6_Result(85) => Dangling_Input_Signal,
       odd6_Result(86) => Dangling_Input_Signal,
       odd6_Result(87) => Dangling_Input_Signal,
       odd6_Result(88) => Dangling_Input_Signal,
       odd6_Result(89) => Dangling_Input_Signal,
       odd6_Result(90) => Dangling_Input_Signal,
       odd6_Result(91) => Dangling_Input_Signal,
       odd6_Result(92) => Dangling_Input_Signal,
       odd6_Result(93) => Dangling_Input_Signal,
       odd6_Result(94) => Dangling_Input_Signal,
       odd6_Result(95) => Dangling_Input_Signal,
       odd6_Result(96) => Dangling_Input_Signal,
       odd6_Result(97) => Dangling_Input_Signal,
       odd6_Result(98) => Dangling_Input_Signal,
       odd6_Result(99) => Dangling_Input_Signal,
       odd6_Result(100) => Dangling_Input_Signal,
       odd6_Result(101) => Dangling_Input_Signal,
       odd6_Result(102) => Dangling_Input_Signal,
       odd6_Result(103) => Dangling_Input_Signal,
       odd6_Result(104) => Dangling_Input_Signal,
       odd6_Result(105) => Dangling_Input_Signal,
       odd6_Result(106) => Dangling_Input_Signal,
       odd6_Result(107) => Dangling_Input_Signal,
       odd6_Result(108) => Dangling_Input_Signal,
       odd6_Result(109) => Dangling_Input_Signal,
       odd6_Result(110) => Dangling_Input_Signal,
       odd6_Result(111) => Dangling_Input_Signal,
       odd6_Result(112) => Dangling_Input_Signal,
       odd6_Result(113) => Dangling_Input_Signal,
       odd6_Result(114) => Dangling_Input_Signal,
       odd6_Result(115) => Dangling_Input_Signal,
       odd6_Result(116) => Dangling_Input_Signal,
       odd6_Result(117) => Dangling_Input_Signal,
       odd6_Result(118) => Dangling_Input_Signal,
       odd6_Result(119) => Dangling_Input_Signal,
       odd6_Result(120) => Dangling_Input_Signal,
       odd6_Result(121) => Dangling_Input_Signal,
       odd6_Result(122) => Dangling_Input_Signal,
       odd6_Result(123) => Dangling_Input_Signal,
       odd6_Result(124) => Dangling_Input_Signal,
       odd6_Result(125) => Dangling_Input_Signal,
       odd6_Result(126) => Dangling_Input_Signal,
       odd6_Result(127) => Dangling_Input_Signal,
       odd7_Latency(0) => Dangling_Input_Signal,
       odd7_Latency(1) => Dangling_Input_Signal,
       odd7_Latency(2) => Dangling_Input_Signal,
       odd7_RegDst(0) => Dangling_Input_Signal,
       odd7_RegDst(1) => Dangling_Input_Signal,
       odd7_RegDst(2) => Dangling_Input_Signal,
       odd7_RegDst(3) => Dangling_Input_Signal,
       odd7_RegDst(4) => Dangling_Input_Signal,
       odd7_RegDst(5) => Dangling_Input_Signal,
       odd7_RegDst(6) => Dangling_Input_Signal,
       odd7_Result(0) => Dangling_Input_Signal,
       odd7_Result(1) => Dangling_Input_Signal,
       odd7_Result(2) => Dangling_Input_Signal,
       odd7_Result(3) => Dangling_Input_Signal,
       odd7_Result(4) => Dangling_Input_Signal,
       odd7_Result(5) => Dangling_Input_Signal,
       odd7_Result(6) => Dangling_Input_Signal,
       odd7_Result(7) => Dangling_Input_Signal,
       odd7_Result(8) => Dangling_Input_Signal,
       odd7_Result(9) => Dangling_Input_Signal,
       odd7_Result(10) => Dangling_Input_Signal,
       odd7_Result(11) => Dangling_Input_Signal,
       odd7_Result(12) => Dangling_Input_Signal,
       odd7_Result(13) => Dangling_Input_Signal,
       odd7_Result(14) => Dangling_Input_Signal,
       odd7_Result(15) => Dangling_Input_Signal,
       odd7_Result(16) => Dangling_Input_Signal,
       odd7_Result(17) => Dangling_Input_Signal,
       odd7_Result(18) => Dangling_Input_Signal,
       odd7_Result(19) => Dangling_Input_Signal,
       odd7_Result(20) => Dangling_Input_Signal,
       odd7_Result(21) => Dangling_Input_Signal,
       odd7_Result(22) => Dangling_Input_Signal,
       odd7_Result(23) => Dangling_Input_Signal,
       odd7_Result(24) => Dangling_Input_Signal,
       odd7_Result(25) => Dangling_Input_Signal,
       odd7_Result(26) => Dangling_Input_Signal,
       odd7_Result(27) => Dangling_Input_Signal,
       odd7_Result(28) => Dangling_Input_Signal,
       odd7_Result(29) => Dangling_Input_Signal,
       odd7_Result(30) => Dangling_Input_Signal,
       odd7_Result(31) => Dangling_Input_Signal,
       odd7_Result(32) => Dangling_Input_Signal,
       odd7_Result(33) => Dangling_Input_Signal,
       odd7_Result(34) => Dangling_Input_Signal,
       odd7_Result(35) => Dangling_Input_Signal,
       odd7_Result(36) => Dangling_Input_Signal,
       odd7_Result(37) => Dangling_Input_Signal,
       odd7_Result(38) => Dangling_Input_Signal,
       odd7_Result(39) => Dangling_Input_Signal,
       odd7_Result(40) => Dangling_Input_Signal,
       odd7_Result(41) => Dangling_Input_Signal,
       odd7_Result(42) => Dangling_Input_Signal,
       odd7_Result(43) => Dangling_Input_Signal,
       odd7_Result(44) => Dangling_Input_Signal,
       odd7_Result(45) => Dangling_Input_Signal,
       odd7_Result(46) => Dangling_Input_Signal,
       odd7_Result(47) => Dangling_Input_Signal,
       odd7_Result(48) => Dangling_Input_Signal,
       odd7_Result(49) => Dangling_Input_Signal,
       odd7_Result(50) => Dangling_Input_Signal,
       odd7_Result(51) => Dangling_Input_Signal,
       odd7_Result(52) => Dangling_Input_Signal,
       odd7_Result(53) => Dangling_Input_Signal,
       odd7_Result(54) => Dangling_Input_Signal,
       odd7_Result(55) => Dangling_Input_Signal,
       odd7_Result(56) => Dangling_Input_Signal,
       odd7_Result(57) => Dangling_Input_Signal,
       odd7_Result(58) => Dangling_Input_Signal,
       odd7_Result(59) => Dangling_Input_Signal,
       odd7_Result(60) => Dangling_Input_Signal,
       odd7_Result(61) => Dangling_Input_Signal,
       odd7_Result(62) => Dangling_Input_Signal,
       odd7_Result(63) => Dangling_Input_Signal,
       odd7_Result(64) => Dangling_Input_Signal,
       odd7_Result(65) => Dangling_Input_Signal,
       odd7_Result(66) => Dangling_Input_Signal,
       odd7_Result(67) => Dangling_Input_Signal,
       odd7_Result(68) => Dangling_Input_Signal,
       odd7_Result(69) => Dangling_Input_Signal,
       odd7_Result(70) => Dangling_Input_Signal,
       odd7_Result(71) => Dangling_Input_Signal,
       odd7_Result(72) => Dangling_Input_Signal,
       odd7_Result(73) => Dangling_Input_Signal,
       odd7_Result(74) => Dangling_Input_Signal,
       odd7_Result(75) => Dangling_Input_Signal,
       odd7_Result(76) => Dangling_Input_Signal,
       odd7_Result(77) => Dangling_Input_Signal,
       odd7_Result(78) => Dangling_Input_Signal,
       odd7_Result(79) => Dangling_Input_Signal,
       odd7_Result(80) => Dangling_Input_Signal,
       odd7_Result(81) => Dangling_Input_Signal,
       odd7_Result(82) => Dangling_Input_Signal,
       odd7_Result(83) => Dangling_Input_Signal,
       odd7_Result(84) => Dangling_Input_Signal,
       odd7_Result(85) => Dangling_Input_Signal,
       odd7_Result(86) => Dangling_Input_Signal,
       odd7_Result(87) => Dangling_Input_Signal,
       odd7_Result(88) => Dangling_Input_Signal,
       odd7_Result(89) => Dangling_Input_Signal,
       odd7_Result(90) => Dangling_Input_Signal,
       odd7_Result(91) => Dangling_Input_Signal,
       odd7_Result(92) => Dangling_Input_Signal,
       odd7_Result(93) => Dangling_Input_Signal,
       odd7_Result(94) => Dangling_Input_Signal,
       odd7_Result(95) => Dangling_Input_Signal,
       odd7_Result(96) => Dangling_Input_Signal,
       odd7_Result(97) => Dangling_Input_Signal,
       odd7_Result(98) => Dangling_Input_Signal,
       odd7_Result(99) => Dangling_Input_Signal,
       odd7_Result(100) => Dangling_Input_Signal,
       odd7_Result(101) => Dangling_Input_Signal,
       odd7_Result(102) => Dangling_Input_Signal,
       odd7_Result(103) => Dangling_Input_Signal,
       odd7_Result(104) => Dangling_Input_Signal,
       odd7_Result(105) => Dangling_Input_Signal,
       odd7_Result(106) => Dangling_Input_Signal,
       odd7_Result(107) => Dangling_Input_Signal,
       odd7_Result(108) => Dangling_Input_Signal,
       odd7_Result(109) => Dangling_Input_Signal,
       odd7_Result(110) => Dangling_Input_Signal,
       odd7_Result(111) => Dangling_Input_Signal,
       odd7_Result(112) => Dangling_Input_Signal,
       odd7_Result(113) => Dangling_Input_Signal,
       odd7_Result(114) => Dangling_Input_Signal,
       odd7_Result(115) => Dangling_Input_Signal,
       odd7_Result(116) => Dangling_Input_Signal,
       odd7_Result(117) => Dangling_Input_Signal,
       odd7_Result(118) => Dangling_Input_Signal,
       odd7_Result(119) => Dangling_Input_Signal,
       odd7_Result(120) => Dangling_Input_Signal,
       odd7_Result(121) => Dangling_Input_Signal,
       odd7_Result(122) => Dangling_Input_Signal,
       odd7_Result(123) => Dangling_Input_Signal,
       odd7_Result(124) => Dangling_Input_Signal,
       odd7_Result(125) => Dangling_Input_Signal,
       odd7_Result(126) => Dangling_Input_Signal,
       odd7_Result(127) => Dangling_Input_Signal,
       RA(0) => Dangling_Input_Signal,
       RA(1) => Dangling_Input_Signal,
       RA(2) => Dangling_Input_Signal,
       RA(3) => Dangling_Input_Signal,
       RA(4) => Dangling_Input_Signal,
       RA(5) => Dangling_Input_Signal,
       RA(6) => Dangling_Input_Signal,
       RB(0) => Dangling_Input_Signal,
       RB(1) => Dangling_Input_Signal,
       RB(2) => Dangling_Input_Signal,
       RB(3) => Dangling_Input_Signal,
       RB(4) => Dangling_Input_Signal,
       RB(5) => Dangling_Input_Signal,
       RB(6) => Dangling_Input_Signal,
       RC(0) => Dangling_Input_Signal,
       RC(1) => Dangling_Input_Signal,
       RC(2) => Dangling_Input_Signal,
       RC(3) => Dangling_Input_Signal,
       RC(4) => Dangling_Input_Signal,
       RC(5) => Dangling_Input_Signal,
       RC(6) => Dangling_Input_Signal,
       RD(0) => Dangling_Input_Signal,
       RD(1) => Dangling_Input_Signal,
       RD(2) => Dangling_Input_Signal,
       RD(3) => Dangling_Input_Signal,
       RD(4) => Dangling_Input_Signal,
       RD(5) => Dangling_Input_Signal,
       RD(6) => Dangling_Input_Signal,
       RE(0) => Dangling_Input_Signal,
       RE(1) => Dangling_Input_Signal,
       RE(2) => Dangling_Input_Signal,
       RE(3) => Dangling_Input_Signal,
       RE(4) => Dangling_Input_Signal,
       RE(5) => Dangling_Input_Signal,
       RE(6) => Dangling_Input_Signal,
       RF(0) => Dangling_Input_Signal,
       RF(1) => Dangling_Input_Signal,
       RF(2) => Dangling_Input_Signal,
       RF(3) => Dangling_Input_Signal,
       RF(4) => Dangling_Input_Signal,
       RF(5) => Dangling_Input_Signal,
       RF(6) => Dangling_Input_Signal,
       even1_RegWr => Dangling_Input_Signal,
       even2_RegWr => Dangling_Input_Signal,
       even3_RegWr => Dangling_Input_Signal,
       even4_RegWr => Dangling_Input_Signal,
       even5_RegWr => Dangling_Input_Signal,
       even6_RegWr => Dangling_Input_Signal,
       even7_RegWr => Dangling_Input_Signal,
       odd1_RegWr => Dangling_Input_Signal,
       odd2_RegWr => Dangling_Input_Signal,
       odd3_RegWr => Dangling_Input_Signal,
       odd4_RegWr => Dangling_Input_Signal,
       odd5_RegWr => Dangling_Input_Signal,
       odd6_RegWr => Dangling_Input_Signal,
       odd7_RegWr => Dangling_Input_Signal
  );


---- Dangling input signal assignment ----

Dangling_Input_Signal <= DANGLING_INPUT_CONSTANT;

end top;
